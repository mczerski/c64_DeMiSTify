
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"d0",x"c8",x"c3",x"87"),
    12 => (x"86",x"c0",x"c6",x"4e"),
    13 => (x"49",x"d0",x"c8",x"c3"),
    14 => (x"48",x"f8",x"f4",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"c3",x"e6"),
    19 => (x"1e",x"87",x"fc",x"98"),
    20 => (x"1e",x"73",x"1e",x"72"),
    21 => (x"02",x"11",x"48",x"12"),
    22 => (x"c3",x"4b",x"87",x"ca"),
    23 => (x"73",x"9b",x"98",x"df"),
    24 => (x"87",x"f0",x"02",x"88"),
    25 => (x"4a",x"26",x"4b",x"26"),
    26 => (x"73",x"1e",x"4f",x"26"),
    27 => (x"c1",x"1e",x"72",x"1e"),
    28 => (x"87",x"ca",x"04",x"8b"),
    29 => (x"02",x"11",x"48",x"12"),
    30 => (x"02",x"88",x"87",x"c4"),
    31 => (x"4a",x"26",x"87",x"f1"),
    32 => (x"4f",x"26",x"4b",x"26"),
    33 => (x"73",x"1e",x"74",x"1e"),
    34 => (x"c1",x"1e",x"72",x"1e"),
    35 => (x"87",x"d0",x"04",x"8b"),
    36 => (x"02",x"11",x"48",x"12"),
    37 => (x"c3",x"4c",x"87",x"ca"),
    38 => (x"74",x"9c",x"98",x"df"),
    39 => (x"87",x"eb",x"02",x"88"),
    40 => (x"4b",x"26",x"4a",x"26"),
    41 => (x"4f",x"26",x"4c",x"26"),
    42 => (x"81",x"48",x"73",x"1e"),
    43 => (x"c5",x"02",x"a9",x"73"),
    44 => (x"05",x"53",x"12",x"87"),
    45 => (x"4f",x"26",x"87",x"f6"),
    46 => (x"4a",x"66",x"c4",x"1e"),
    47 => (x"51",x"12",x"48",x"71"),
    48 => (x"26",x"87",x"fb",x"05"),
    49 => (x"4a",x"71",x"1e",x"4f"),
    50 => (x"48",x"49",x"66",x"c4"),
    51 => (x"a6",x"c8",x"88",x"c1"),
    52 => (x"02",x"99",x"71",x"58"),
    53 => (x"48",x"12",x"87",x"d4"),
    54 => (x"78",x"08",x"d4",x"ff"),
    55 => (x"48",x"49",x"66",x"c4"),
    56 => (x"a6",x"c8",x"88",x"c1"),
    57 => (x"05",x"99",x"71",x"58"),
    58 => (x"4f",x"26",x"87",x"ec"),
    59 => (x"c4",x"4a",x"71",x"1e"),
    60 => (x"c1",x"48",x"49",x"66"),
    61 => (x"58",x"a6",x"c8",x"88"),
    62 => (x"d6",x"02",x"99",x"71"),
    63 => (x"48",x"d4",x"ff",x"87"),
    64 => (x"68",x"78",x"ff",x"c3"),
    65 => (x"49",x"66",x"c4",x"52"),
    66 => (x"c8",x"88",x"c1",x"48"),
    67 => (x"99",x"71",x"58",x"a6"),
    68 => (x"26",x"87",x"ea",x"05"),
    69 => (x"1e",x"73",x"1e",x"4f"),
    70 => (x"c3",x"4b",x"d4",x"ff"),
    71 => (x"4a",x"6b",x"7b",x"ff"),
    72 => (x"6b",x"7b",x"ff",x"c3"),
    73 => (x"72",x"32",x"c8",x"49"),
    74 => (x"7b",x"ff",x"c3",x"b1"),
    75 => (x"31",x"c8",x"4a",x"6b"),
    76 => (x"ff",x"c3",x"b2",x"71"),
    77 => (x"c8",x"49",x"6b",x"7b"),
    78 => (x"71",x"b1",x"72",x"32"),
    79 => (x"26",x"87",x"c4",x"48"),
    80 => (x"26",x"4c",x"26",x"4d"),
    81 => (x"0e",x"4f",x"26",x"4b"),
    82 => (x"5d",x"5c",x"5b",x"5e"),
    83 => (x"ff",x"4a",x"71",x"0e"),
    84 => (x"49",x"72",x"4c",x"d4"),
    85 => (x"71",x"99",x"ff",x"c3"),
    86 => (x"f8",x"f4",x"c2",x"7c"),
    87 => (x"87",x"c8",x"05",x"bf"),
    88 => (x"c9",x"48",x"66",x"d0"),
    89 => (x"58",x"a6",x"d4",x"30"),
    90 => (x"d8",x"49",x"66",x"d0"),
    91 => (x"99",x"ff",x"c3",x"29"),
    92 => (x"66",x"d0",x"7c",x"71"),
    93 => (x"c3",x"29",x"d0",x"49"),
    94 => (x"7c",x"71",x"99",x"ff"),
    95 => (x"c8",x"49",x"66",x"d0"),
    96 => (x"99",x"ff",x"c3",x"29"),
    97 => (x"66",x"d0",x"7c",x"71"),
    98 => (x"99",x"ff",x"c3",x"49"),
    99 => (x"49",x"72",x"7c",x"71"),
   100 => (x"ff",x"c3",x"29",x"d0"),
   101 => (x"6c",x"7c",x"71",x"99"),
   102 => (x"ff",x"f0",x"c9",x"4b"),
   103 => (x"ab",x"ff",x"c3",x"4d"),
   104 => (x"c3",x"87",x"d0",x"05"),
   105 => (x"4b",x"6c",x"7c",x"ff"),
   106 => (x"c6",x"02",x"8d",x"c1"),
   107 => (x"ab",x"ff",x"c3",x"87"),
   108 => (x"73",x"87",x"f0",x"02"),
   109 => (x"87",x"c7",x"fe",x"48"),
   110 => (x"ff",x"49",x"c0",x"1e"),
   111 => (x"ff",x"c3",x"48",x"d4"),
   112 => (x"c3",x"81",x"c1",x"78"),
   113 => (x"04",x"a9",x"b7",x"c8"),
   114 => (x"4f",x"26",x"87",x"f1"),
   115 => (x"e7",x"1e",x"73",x"1e"),
   116 => (x"df",x"f8",x"c4",x"87"),
   117 => (x"c0",x"1e",x"c0",x"4b"),
   118 => (x"f7",x"c1",x"f0",x"ff"),
   119 => (x"87",x"e7",x"fd",x"49"),
   120 => (x"a8",x"c1",x"86",x"c4"),
   121 => (x"87",x"ea",x"c0",x"05"),
   122 => (x"c3",x"48",x"d4",x"ff"),
   123 => (x"c0",x"c1",x"78",x"ff"),
   124 => (x"c0",x"c0",x"c0",x"c0"),
   125 => (x"f0",x"e1",x"c0",x"1e"),
   126 => (x"fd",x"49",x"e9",x"c1"),
   127 => (x"86",x"c4",x"87",x"c9"),
   128 => (x"ca",x"05",x"98",x"70"),
   129 => (x"48",x"d4",x"ff",x"87"),
   130 => (x"c1",x"78",x"ff",x"c3"),
   131 => (x"fe",x"87",x"cb",x"48"),
   132 => (x"8b",x"c1",x"87",x"e6"),
   133 => (x"87",x"fd",x"fe",x"05"),
   134 => (x"e6",x"fc",x"48",x"c0"),
   135 => (x"1e",x"73",x"1e",x"87"),
   136 => (x"c3",x"48",x"d4",x"ff"),
   137 => (x"4b",x"d3",x"78",x"ff"),
   138 => (x"ff",x"c0",x"1e",x"c0"),
   139 => (x"49",x"c1",x"c1",x"f0"),
   140 => (x"c4",x"87",x"d4",x"fc"),
   141 => (x"05",x"98",x"70",x"86"),
   142 => (x"d4",x"ff",x"87",x"ca"),
   143 => (x"78",x"ff",x"c3",x"48"),
   144 => (x"87",x"cb",x"48",x"c1"),
   145 => (x"c1",x"87",x"f1",x"fd"),
   146 => (x"db",x"ff",x"05",x"8b"),
   147 => (x"fb",x"48",x"c0",x"87"),
   148 => (x"5e",x"0e",x"87",x"f1"),
   149 => (x"ff",x"0e",x"5c",x"5b"),
   150 => (x"db",x"fd",x"4c",x"d4"),
   151 => (x"1e",x"ea",x"c6",x"87"),
   152 => (x"c1",x"f0",x"e1",x"c0"),
   153 => (x"de",x"fb",x"49",x"c8"),
   154 => (x"c1",x"86",x"c4",x"87"),
   155 => (x"87",x"c8",x"02",x"a8"),
   156 => (x"c0",x"87",x"ea",x"fe"),
   157 => (x"87",x"e2",x"c1",x"48"),
   158 => (x"70",x"87",x"da",x"fa"),
   159 => (x"ff",x"ff",x"cf",x"49"),
   160 => (x"a9",x"ea",x"c6",x"99"),
   161 => (x"fe",x"87",x"c8",x"02"),
   162 => (x"48",x"c0",x"87",x"d3"),
   163 => (x"c3",x"87",x"cb",x"c1"),
   164 => (x"f1",x"c0",x"7c",x"ff"),
   165 => (x"87",x"f4",x"fc",x"4b"),
   166 => (x"c0",x"02",x"98",x"70"),
   167 => (x"1e",x"c0",x"87",x"eb"),
   168 => (x"c1",x"f0",x"ff",x"c0"),
   169 => (x"de",x"fa",x"49",x"fa"),
   170 => (x"70",x"86",x"c4",x"87"),
   171 => (x"87",x"d9",x"05",x"98"),
   172 => (x"6c",x"7c",x"ff",x"c3"),
   173 => (x"7c",x"ff",x"c3",x"49"),
   174 => (x"c1",x"7c",x"7c",x"7c"),
   175 => (x"c4",x"02",x"99",x"c0"),
   176 => (x"d5",x"48",x"c1",x"87"),
   177 => (x"d1",x"48",x"c0",x"87"),
   178 => (x"05",x"ab",x"c2",x"87"),
   179 => (x"48",x"c0",x"87",x"c4"),
   180 => (x"8b",x"c1",x"87",x"c8"),
   181 => (x"87",x"fd",x"fe",x"05"),
   182 => (x"e4",x"f9",x"48",x"c0"),
   183 => (x"1e",x"73",x"1e",x"87"),
   184 => (x"48",x"f8",x"f4",x"c2"),
   185 => (x"4b",x"c7",x"78",x"c1"),
   186 => (x"c2",x"48",x"d0",x"ff"),
   187 => (x"87",x"c8",x"fb",x"78"),
   188 => (x"c3",x"48",x"d0",x"ff"),
   189 => (x"c0",x"1e",x"c0",x"78"),
   190 => (x"c0",x"c1",x"d0",x"e5"),
   191 => (x"87",x"c7",x"f9",x"49"),
   192 => (x"a8",x"c1",x"86",x"c4"),
   193 => (x"4b",x"87",x"c1",x"05"),
   194 => (x"c5",x"05",x"ab",x"c2"),
   195 => (x"c0",x"48",x"c0",x"87"),
   196 => (x"8b",x"c1",x"87",x"f9"),
   197 => (x"87",x"d0",x"ff",x"05"),
   198 => (x"c2",x"87",x"f7",x"fc"),
   199 => (x"70",x"58",x"fc",x"f4"),
   200 => (x"87",x"cd",x"05",x"98"),
   201 => (x"ff",x"c0",x"1e",x"c1"),
   202 => (x"49",x"d0",x"c1",x"f0"),
   203 => (x"c4",x"87",x"d8",x"f8"),
   204 => (x"48",x"d4",x"ff",x"86"),
   205 => (x"c4",x"78",x"ff",x"c3"),
   206 => (x"f5",x"c2",x"87",x"de"),
   207 => (x"d0",x"ff",x"58",x"c0"),
   208 => (x"ff",x"78",x"c2",x"48"),
   209 => (x"ff",x"c3",x"48",x"d4"),
   210 => (x"f7",x"48",x"c1",x"78"),
   211 => (x"5e",x"0e",x"87",x"f5"),
   212 => (x"0e",x"5d",x"5c",x"5b"),
   213 => (x"ff",x"c3",x"4a",x"71"),
   214 => (x"4c",x"d4",x"ff",x"4d"),
   215 => (x"d0",x"ff",x"7c",x"75"),
   216 => (x"78",x"c3",x"c4",x"48"),
   217 => (x"1e",x"72",x"7c",x"75"),
   218 => (x"c1",x"f0",x"ff",x"c0"),
   219 => (x"d6",x"f7",x"49",x"d8"),
   220 => (x"70",x"86",x"c4",x"87"),
   221 => (x"87",x"c5",x"02",x"98"),
   222 => (x"f0",x"c0",x"48",x"c1"),
   223 => (x"c3",x"7c",x"75",x"87"),
   224 => (x"c0",x"c8",x"7c",x"fe"),
   225 => (x"49",x"66",x"d4",x"1e"),
   226 => (x"c4",x"87",x"fa",x"f4"),
   227 => (x"75",x"7c",x"75",x"86"),
   228 => (x"d8",x"7c",x"75",x"7c"),
   229 => (x"75",x"4b",x"e0",x"da"),
   230 => (x"99",x"49",x"6c",x"7c"),
   231 => (x"c1",x"87",x"c5",x"05"),
   232 => (x"87",x"f3",x"05",x"8b"),
   233 => (x"d0",x"ff",x"7c",x"75"),
   234 => (x"c0",x"78",x"c2",x"48"),
   235 => (x"87",x"cf",x"f6",x"48"),
   236 => (x"5c",x"5b",x"5e",x"0e"),
   237 => (x"4b",x"71",x"0e",x"5d"),
   238 => (x"ee",x"c5",x"4c",x"c0"),
   239 => (x"ff",x"4a",x"df",x"cd"),
   240 => (x"ff",x"c3",x"48",x"d4"),
   241 => (x"c3",x"49",x"68",x"78"),
   242 => (x"c0",x"05",x"a9",x"fe"),
   243 => (x"4d",x"70",x"87",x"fd"),
   244 => (x"cc",x"02",x"9b",x"73"),
   245 => (x"1e",x"66",x"d0",x"87"),
   246 => (x"cf",x"f4",x"49",x"73"),
   247 => (x"d6",x"86",x"c4",x"87"),
   248 => (x"48",x"d0",x"ff",x"87"),
   249 => (x"c3",x"78",x"d1",x"c4"),
   250 => (x"66",x"d0",x"7d",x"ff"),
   251 => (x"d4",x"88",x"c1",x"48"),
   252 => (x"98",x"70",x"58",x"a6"),
   253 => (x"ff",x"87",x"f0",x"05"),
   254 => (x"ff",x"c3",x"48",x"d4"),
   255 => (x"9b",x"73",x"78",x"78"),
   256 => (x"ff",x"87",x"c5",x"05"),
   257 => (x"78",x"d0",x"48",x"d0"),
   258 => (x"c1",x"4c",x"4a",x"c1"),
   259 => (x"ee",x"fe",x"05",x"8a"),
   260 => (x"f4",x"48",x"74",x"87"),
   261 => (x"73",x"1e",x"87",x"e9"),
   262 => (x"c0",x"4a",x"71",x"1e"),
   263 => (x"48",x"d4",x"ff",x"4b"),
   264 => (x"ff",x"78",x"ff",x"c3"),
   265 => (x"c3",x"c4",x"48",x"d0"),
   266 => (x"48",x"d4",x"ff",x"78"),
   267 => (x"72",x"78",x"ff",x"c3"),
   268 => (x"f0",x"ff",x"c0",x"1e"),
   269 => (x"f4",x"49",x"d1",x"c1"),
   270 => (x"86",x"c4",x"87",x"cd"),
   271 => (x"d2",x"05",x"98",x"70"),
   272 => (x"1e",x"c0",x"c8",x"87"),
   273 => (x"fd",x"49",x"66",x"cc"),
   274 => (x"86",x"c4",x"87",x"e6"),
   275 => (x"d0",x"ff",x"4b",x"70"),
   276 => (x"73",x"78",x"c2",x"48"),
   277 => (x"87",x"eb",x"f3",x"48"),
   278 => (x"5c",x"5b",x"5e",x"0e"),
   279 => (x"1e",x"c0",x"0e",x"5d"),
   280 => (x"c1",x"f0",x"ff",x"c0"),
   281 => (x"de",x"f3",x"49",x"c9"),
   282 => (x"c2",x"1e",x"d2",x"87"),
   283 => (x"fc",x"49",x"c0",x"f5"),
   284 => (x"86",x"c8",x"87",x"fe"),
   285 => (x"84",x"c1",x"4c",x"c0"),
   286 => (x"04",x"ac",x"b7",x"d2"),
   287 => (x"f5",x"c2",x"87",x"f8"),
   288 => (x"49",x"bf",x"97",x"c0"),
   289 => (x"c1",x"99",x"c0",x"c3"),
   290 => (x"c0",x"05",x"a9",x"c0"),
   291 => (x"f5",x"c2",x"87",x"e7"),
   292 => (x"49",x"bf",x"97",x"c7"),
   293 => (x"f5",x"c2",x"31",x"d0"),
   294 => (x"4a",x"bf",x"97",x"c8"),
   295 => (x"b1",x"72",x"32",x"c8"),
   296 => (x"97",x"c9",x"f5",x"c2"),
   297 => (x"71",x"b1",x"4a",x"bf"),
   298 => (x"ff",x"ff",x"cf",x"4c"),
   299 => (x"84",x"c1",x"9c",x"ff"),
   300 => (x"e7",x"c1",x"34",x"ca"),
   301 => (x"c9",x"f5",x"c2",x"87"),
   302 => (x"c1",x"49",x"bf",x"97"),
   303 => (x"c2",x"99",x"c6",x"31"),
   304 => (x"bf",x"97",x"ca",x"f5"),
   305 => (x"2a",x"b7",x"c7",x"4a"),
   306 => (x"f5",x"c2",x"b1",x"72"),
   307 => (x"4a",x"bf",x"97",x"c5"),
   308 => (x"c2",x"9d",x"cf",x"4d"),
   309 => (x"bf",x"97",x"c6",x"f5"),
   310 => (x"ca",x"9a",x"c3",x"4a"),
   311 => (x"c7",x"f5",x"c2",x"32"),
   312 => (x"c2",x"4b",x"bf",x"97"),
   313 => (x"c2",x"b2",x"73",x"33"),
   314 => (x"bf",x"97",x"c8",x"f5"),
   315 => (x"9b",x"c0",x"c3",x"4b"),
   316 => (x"73",x"2b",x"b7",x"c6"),
   317 => (x"c1",x"81",x"c2",x"b2"),
   318 => (x"70",x"30",x"71",x"48"),
   319 => (x"75",x"48",x"c1",x"49"),
   320 => (x"72",x"4d",x"70",x"30"),
   321 => (x"71",x"84",x"c1",x"4c"),
   322 => (x"b7",x"c0",x"c8",x"94"),
   323 => (x"87",x"cc",x"06",x"ad"),
   324 => (x"2d",x"b7",x"34",x"c1"),
   325 => (x"ad",x"b7",x"c0",x"c8"),
   326 => (x"87",x"f4",x"ff",x"01"),
   327 => (x"de",x"f0",x"48",x"74"),
   328 => (x"5b",x"5e",x"0e",x"87"),
   329 => (x"f8",x"0e",x"5d",x"5c"),
   330 => (x"e6",x"fd",x"c2",x"86"),
   331 => (x"c2",x"78",x"c0",x"48"),
   332 => (x"c0",x"1e",x"de",x"f5"),
   333 => (x"87",x"de",x"fb",x"49"),
   334 => (x"98",x"70",x"86",x"c4"),
   335 => (x"c0",x"87",x"c5",x"05"),
   336 => (x"87",x"ce",x"c9",x"48"),
   337 => (x"7e",x"c1",x"4d",x"c0"),
   338 => (x"bf",x"c0",x"f3",x"c0"),
   339 => (x"d4",x"f6",x"c2",x"49"),
   340 => (x"4b",x"c8",x"71",x"4a"),
   341 => (x"70",x"87",x"d3",x"ec"),
   342 => (x"87",x"c2",x"05",x"98"),
   343 => (x"f2",x"c0",x"7e",x"c0"),
   344 => (x"c2",x"49",x"bf",x"fc"),
   345 => (x"71",x"4a",x"f0",x"f6"),
   346 => (x"fd",x"eb",x"4b",x"c8"),
   347 => (x"05",x"98",x"70",x"87"),
   348 => (x"7e",x"c0",x"87",x"c2"),
   349 => (x"fd",x"c0",x"02",x"6e"),
   350 => (x"e4",x"fc",x"c2",x"87"),
   351 => (x"fd",x"c2",x"4d",x"bf"),
   352 => (x"7e",x"bf",x"9f",x"dc"),
   353 => (x"ea",x"d6",x"c5",x"48"),
   354 => (x"87",x"c7",x"05",x"a8"),
   355 => (x"bf",x"e4",x"fc",x"c2"),
   356 => (x"6e",x"87",x"ce",x"4d"),
   357 => (x"d5",x"e9",x"ca",x"48"),
   358 => (x"87",x"c5",x"02",x"a8"),
   359 => (x"f1",x"c7",x"48",x"c0"),
   360 => (x"de",x"f5",x"c2",x"87"),
   361 => (x"f9",x"49",x"75",x"1e"),
   362 => (x"86",x"c4",x"87",x"ec"),
   363 => (x"c5",x"05",x"98",x"70"),
   364 => (x"c7",x"48",x"c0",x"87"),
   365 => (x"f2",x"c0",x"87",x"dc"),
   366 => (x"c2",x"49",x"bf",x"fc"),
   367 => (x"71",x"4a",x"f0",x"f6"),
   368 => (x"e5",x"ea",x"4b",x"c8"),
   369 => (x"05",x"98",x"70",x"87"),
   370 => (x"fd",x"c2",x"87",x"c8"),
   371 => (x"78",x"c1",x"48",x"e6"),
   372 => (x"f3",x"c0",x"87",x"da"),
   373 => (x"c2",x"49",x"bf",x"c0"),
   374 => (x"71",x"4a",x"d4",x"f6"),
   375 => (x"c9",x"ea",x"4b",x"c8"),
   376 => (x"02",x"98",x"70",x"87"),
   377 => (x"c0",x"87",x"c5",x"c0"),
   378 => (x"87",x"e6",x"c6",x"48"),
   379 => (x"97",x"dc",x"fd",x"c2"),
   380 => (x"d5",x"c1",x"49",x"bf"),
   381 => (x"cd",x"c0",x"05",x"a9"),
   382 => (x"dd",x"fd",x"c2",x"87"),
   383 => (x"c2",x"49",x"bf",x"97"),
   384 => (x"c0",x"02",x"a9",x"ea"),
   385 => (x"48",x"c0",x"87",x"c5"),
   386 => (x"c2",x"87",x"c7",x"c6"),
   387 => (x"bf",x"97",x"de",x"f5"),
   388 => (x"e9",x"c3",x"48",x"7e"),
   389 => (x"ce",x"c0",x"02",x"a8"),
   390 => (x"c3",x"48",x"6e",x"87"),
   391 => (x"c0",x"02",x"a8",x"eb"),
   392 => (x"48",x"c0",x"87",x"c5"),
   393 => (x"c2",x"87",x"eb",x"c5"),
   394 => (x"bf",x"97",x"e9",x"f5"),
   395 => (x"c0",x"05",x"99",x"49"),
   396 => (x"f5",x"c2",x"87",x"cc"),
   397 => (x"49",x"bf",x"97",x"ea"),
   398 => (x"c0",x"02",x"a9",x"c2"),
   399 => (x"48",x"c0",x"87",x"c5"),
   400 => (x"c2",x"87",x"cf",x"c5"),
   401 => (x"bf",x"97",x"eb",x"f5"),
   402 => (x"e2",x"fd",x"c2",x"48"),
   403 => (x"48",x"4c",x"70",x"58"),
   404 => (x"fd",x"c2",x"88",x"c1"),
   405 => (x"f5",x"c2",x"58",x"e6"),
   406 => (x"49",x"bf",x"97",x"ec"),
   407 => (x"f5",x"c2",x"81",x"75"),
   408 => (x"4a",x"bf",x"97",x"ed"),
   409 => (x"a1",x"72",x"32",x"c8"),
   410 => (x"f3",x"c1",x"c3",x"7e"),
   411 => (x"c2",x"78",x"6e",x"48"),
   412 => (x"bf",x"97",x"ee",x"f5"),
   413 => (x"58",x"a6",x"c8",x"48"),
   414 => (x"bf",x"e6",x"fd",x"c2"),
   415 => (x"87",x"d4",x"c2",x"02"),
   416 => (x"bf",x"fc",x"f2",x"c0"),
   417 => (x"f0",x"f6",x"c2",x"49"),
   418 => (x"4b",x"c8",x"71",x"4a"),
   419 => (x"70",x"87",x"db",x"e7"),
   420 => (x"c5",x"c0",x"02",x"98"),
   421 => (x"c3",x"48",x"c0",x"87"),
   422 => (x"fd",x"c2",x"87",x"f8"),
   423 => (x"c3",x"4c",x"bf",x"de"),
   424 => (x"c2",x"5c",x"c7",x"c2"),
   425 => (x"bf",x"97",x"c3",x"f6"),
   426 => (x"c2",x"31",x"c8",x"49"),
   427 => (x"bf",x"97",x"c2",x"f6"),
   428 => (x"c2",x"49",x"a1",x"4a"),
   429 => (x"bf",x"97",x"c4",x"f6"),
   430 => (x"72",x"32",x"d0",x"4a"),
   431 => (x"f6",x"c2",x"49",x"a1"),
   432 => (x"4a",x"bf",x"97",x"c5"),
   433 => (x"a1",x"72",x"32",x"d8"),
   434 => (x"91",x"66",x"c4",x"49"),
   435 => (x"bf",x"f3",x"c1",x"c3"),
   436 => (x"fb",x"c1",x"c3",x"81"),
   437 => (x"cb",x"f6",x"c2",x"59"),
   438 => (x"c8",x"4a",x"bf",x"97"),
   439 => (x"ca",x"f6",x"c2",x"32"),
   440 => (x"a2",x"4b",x"bf",x"97"),
   441 => (x"cc",x"f6",x"c2",x"4a"),
   442 => (x"d0",x"4b",x"bf",x"97"),
   443 => (x"4a",x"a2",x"73",x"33"),
   444 => (x"97",x"cd",x"f6",x"c2"),
   445 => (x"9b",x"cf",x"4b",x"bf"),
   446 => (x"a2",x"73",x"33",x"d8"),
   447 => (x"ff",x"c1",x"c3",x"4a"),
   448 => (x"fb",x"c1",x"c3",x"5a"),
   449 => (x"8a",x"c2",x"4a",x"bf"),
   450 => (x"c1",x"c3",x"92",x"74"),
   451 => (x"a1",x"72",x"48",x"ff"),
   452 => (x"87",x"ca",x"c1",x"78"),
   453 => (x"97",x"f0",x"f5",x"c2"),
   454 => (x"31",x"c8",x"49",x"bf"),
   455 => (x"97",x"ef",x"f5",x"c2"),
   456 => (x"49",x"a1",x"4a",x"bf"),
   457 => (x"59",x"ee",x"fd",x"c2"),
   458 => (x"bf",x"ea",x"fd",x"c2"),
   459 => (x"c7",x"31",x"c5",x"49"),
   460 => (x"29",x"c9",x"81",x"ff"),
   461 => (x"59",x"c7",x"c2",x"c3"),
   462 => (x"97",x"f5",x"f5",x"c2"),
   463 => (x"32",x"c8",x"4a",x"bf"),
   464 => (x"97",x"f4",x"f5",x"c2"),
   465 => (x"4a",x"a2",x"4b",x"bf"),
   466 => (x"6e",x"92",x"66",x"c4"),
   467 => (x"c3",x"c2",x"c3",x"82"),
   468 => (x"fb",x"c1",x"c3",x"5a"),
   469 => (x"c3",x"78",x"c0",x"48"),
   470 => (x"72",x"48",x"f7",x"c1"),
   471 => (x"c2",x"c3",x"78",x"a1"),
   472 => (x"c1",x"c3",x"48",x"c7"),
   473 => (x"c3",x"78",x"bf",x"fb"),
   474 => (x"c3",x"48",x"cb",x"c2"),
   475 => (x"78",x"bf",x"ff",x"c1"),
   476 => (x"bf",x"e6",x"fd",x"c2"),
   477 => (x"87",x"c9",x"c0",x"02"),
   478 => (x"30",x"c4",x"48",x"74"),
   479 => (x"c9",x"c0",x"7e",x"70"),
   480 => (x"c3",x"c2",x"c3",x"87"),
   481 => (x"30",x"c4",x"48",x"bf"),
   482 => (x"fd",x"c2",x"7e",x"70"),
   483 => (x"78",x"6e",x"48",x"ea"),
   484 => (x"8e",x"f8",x"48",x"c1"),
   485 => (x"4c",x"26",x"4d",x"26"),
   486 => (x"4f",x"26",x"4b",x"26"),
   487 => (x"5c",x"5b",x"5e",x"0e"),
   488 => (x"4a",x"71",x"0e",x"5d"),
   489 => (x"bf",x"e6",x"fd",x"c2"),
   490 => (x"72",x"87",x"cb",x"02"),
   491 => (x"72",x"2b",x"c7",x"4b"),
   492 => (x"9c",x"ff",x"c1",x"4c"),
   493 => (x"4b",x"72",x"87",x"c9"),
   494 => (x"4c",x"72",x"2b",x"c8"),
   495 => (x"c3",x"9c",x"ff",x"c3"),
   496 => (x"83",x"bf",x"f3",x"c1"),
   497 => (x"bf",x"f8",x"f2",x"c0"),
   498 => (x"87",x"d9",x"02",x"ab"),
   499 => (x"5b",x"fc",x"f2",x"c0"),
   500 => (x"1e",x"de",x"f5",x"c2"),
   501 => (x"fd",x"f0",x"49",x"73"),
   502 => (x"70",x"86",x"c4",x"87"),
   503 => (x"87",x"c5",x"05",x"98"),
   504 => (x"e6",x"c0",x"48",x"c0"),
   505 => (x"e6",x"fd",x"c2",x"87"),
   506 => (x"87",x"d2",x"02",x"bf"),
   507 => (x"91",x"c4",x"49",x"74"),
   508 => (x"81",x"de",x"f5",x"c2"),
   509 => (x"ff",x"cf",x"4d",x"69"),
   510 => (x"9d",x"ff",x"ff",x"ff"),
   511 => (x"49",x"74",x"87",x"cb"),
   512 => (x"f5",x"c2",x"91",x"c2"),
   513 => (x"69",x"9f",x"81",x"de"),
   514 => (x"fe",x"48",x"75",x"4d"),
   515 => (x"5e",x"0e",x"87",x"c6"),
   516 => (x"0e",x"5d",x"5c",x"5b"),
   517 => (x"c0",x"4d",x"71",x"1e"),
   518 => (x"ca",x"49",x"c1",x"1e"),
   519 => (x"86",x"c4",x"87",x"ff"),
   520 => (x"02",x"9c",x"4c",x"70"),
   521 => (x"c2",x"87",x"c0",x"c1"),
   522 => (x"75",x"4a",x"ee",x"fd"),
   523 => (x"87",x"df",x"e0",x"49"),
   524 => (x"c0",x"02",x"98",x"70"),
   525 => (x"4a",x"74",x"87",x"f1"),
   526 => (x"4b",x"cb",x"49",x"75"),
   527 => (x"70",x"87",x"c5",x"e1"),
   528 => (x"e2",x"c0",x"02",x"98"),
   529 => (x"74",x"1e",x"c0",x"87"),
   530 => (x"87",x"c7",x"02",x"9c"),
   531 => (x"c0",x"48",x"a6",x"c4"),
   532 => (x"c4",x"87",x"c5",x"78"),
   533 => (x"78",x"c1",x"48",x"a6"),
   534 => (x"c9",x"49",x"66",x"c4"),
   535 => (x"86",x"c4",x"87",x"ff"),
   536 => (x"05",x"9c",x"4c",x"70"),
   537 => (x"74",x"87",x"c0",x"ff"),
   538 => (x"e7",x"fc",x"26",x"48"),
   539 => (x"5b",x"5e",x"0e",x"87"),
   540 => (x"1e",x"0e",x"5d",x"5c"),
   541 => (x"05",x"9b",x"4b",x"71"),
   542 => (x"48",x"c0",x"87",x"c5"),
   543 => (x"c8",x"87",x"e5",x"c1"),
   544 => (x"7d",x"c0",x"4d",x"a3"),
   545 => (x"c7",x"02",x"66",x"d4"),
   546 => (x"97",x"66",x"d4",x"87"),
   547 => (x"87",x"c5",x"05",x"bf"),
   548 => (x"cf",x"c1",x"48",x"c0"),
   549 => (x"49",x"66",x"d4",x"87"),
   550 => (x"70",x"87",x"f3",x"fd"),
   551 => (x"c1",x"02",x"9c",x"4c"),
   552 => (x"a4",x"dc",x"87",x"c0"),
   553 => (x"da",x"7d",x"69",x"49"),
   554 => (x"a3",x"c4",x"49",x"a4"),
   555 => (x"7a",x"69",x"9f",x"4a"),
   556 => (x"bf",x"e6",x"fd",x"c2"),
   557 => (x"d4",x"87",x"d2",x"02"),
   558 => (x"69",x"9f",x"49",x"a4"),
   559 => (x"ff",x"ff",x"c0",x"49"),
   560 => (x"d0",x"48",x"71",x"99"),
   561 => (x"c2",x"7e",x"70",x"30"),
   562 => (x"6e",x"7e",x"c0",x"87"),
   563 => (x"80",x"6a",x"48",x"49"),
   564 => (x"7b",x"c0",x"7a",x"70"),
   565 => (x"6a",x"49",x"a3",x"cc"),
   566 => (x"49",x"a3",x"d0",x"79"),
   567 => (x"48",x"c1",x"79",x"c0"),
   568 => (x"48",x"c0",x"87",x"c2"),
   569 => (x"87",x"ec",x"fa",x"26"),
   570 => (x"5c",x"5b",x"5e",x"0e"),
   571 => (x"4c",x"71",x"0e",x"5d"),
   572 => (x"ca",x"c1",x"02",x"9c"),
   573 => (x"49",x"a4",x"c8",x"87"),
   574 => (x"c2",x"c1",x"02",x"69"),
   575 => (x"4a",x"66",x"d0",x"87"),
   576 => (x"d4",x"82",x"49",x"6c"),
   577 => (x"66",x"d0",x"5a",x"a6"),
   578 => (x"fd",x"c2",x"b9",x"4d"),
   579 => (x"ff",x"4a",x"bf",x"e2"),
   580 => (x"71",x"99",x"72",x"ba"),
   581 => (x"e4",x"c0",x"02",x"99"),
   582 => (x"4b",x"a4",x"c4",x"87"),
   583 => (x"fb",x"f9",x"49",x"6b"),
   584 => (x"c2",x"7b",x"70",x"87"),
   585 => (x"49",x"bf",x"de",x"fd"),
   586 => (x"7c",x"71",x"81",x"6c"),
   587 => (x"fd",x"c2",x"b9",x"75"),
   588 => (x"ff",x"4a",x"bf",x"e2"),
   589 => (x"71",x"99",x"72",x"ba"),
   590 => (x"dc",x"ff",x"05",x"99"),
   591 => (x"f9",x"7c",x"75",x"87"),
   592 => (x"73",x"1e",x"87",x"d2"),
   593 => (x"9b",x"4b",x"71",x"1e"),
   594 => (x"c8",x"87",x"c7",x"02"),
   595 => (x"05",x"69",x"49",x"a3"),
   596 => (x"48",x"c0",x"87",x"c5"),
   597 => (x"c3",x"87",x"f7",x"c0"),
   598 => (x"4a",x"bf",x"f7",x"c1"),
   599 => (x"69",x"49",x"a3",x"c4"),
   600 => (x"c2",x"89",x"c2",x"49"),
   601 => (x"91",x"bf",x"de",x"fd"),
   602 => (x"c2",x"4a",x"a2",x"71"),
   603 => (x"49",x"bf",x"e2",x"fd"),
   604 => (x"a2",x"71",x"99",x"6b"),
   605 => (x"fc",x"f2",x"c0",x"4a"),
   606 => (x"1e",x"66",x"c8",x"5a"),
   607 => (x"d5",x"ea",x"49",x"72"),
   608 => (x"70",x"86",x"c4",x"87"),
   609 => (x"87",x"c4",x"05",x"98"),
   610 => (x"87",x"c2",x"48",x"c0"),
   611 => (x"c7",x"f8",x"48",x"c1"),
   612 => (x"1e",x"73",x"1e",x"87"),
   613 => (x"02",x"9b",x"4b",x"71"),
   614 => (x"a3",x"c8",x"87",x"c7"),
   615 => (x"c5",x"05",x"69",x"49"),
   616 => (x"c0",x"48",x"c0",x"87"),
   617 => (x"c1",x"c3",x"87",x"f7"),
   618 => (x"c4",x"4a",x"bf",x"f7"),
   619 => (x"49",x"69",x"49",x"a3"),
   620 => (x"fd",x"c2",x"89",x"c2"),
   621 => (x"71",x"91",x"bf",x"de"),
   622 => (x"fd",x"c2",x"4a",x"a2"),
   623 => (x"6b",x"49",x"bf",x"e2"),
   624 => (x"4a",x"a2",x"71",x"99"),
   625 => (x"5a",x"fc",x"f2",x"c0"),
   626 => (x"72",x"1e",x"66",x"c8"),
   627 => (x"87",x"fe",x"e5",x"49"),
   628 => (x"98",x"70",x"86",x"c4"),
   629 => (x"c0",x"87",x"c4",x"05"),
   630 => (x"c1",x"87",x"c2",x"48"),
   631 => (x"87",x"f8",x"f6",x"48"),
   632 => (x"5c",x"5b",x"5e",x"0e"),
   633 => (x"71",x"1e",x"0e",x"5d"),
   634 => (x"4c",x"66",x"d4",x"4b"),
   635 => (x"9b",x"73",x"2c",x"c9"),
   636 => (x"87",x"cf",x"c1",x"02"),
   637 => (x"69",x"49",x"a3",x"c8"),
   638 => (x"87",x"c7",x"c1",x"02"),
   639 => (x"d4",x"4d",x"a3",x"d0"),
   640 => (x"fd",x"c2",x"7d",x"66"),
   641 => (x"ff",x"49",x"bf",x"e2"),
   642 => (x"99",x"4a",x"6b",x"b9"),
   643 => (x"03",x"ac",x"71",x"7e"),
   644 => (x"7b",x"c0",x"87",x"cd"),
   645 => (x"4a",x"a3",x"cc",x"7d"),
   646 => (x"6a",x"49",x"a3",x"c4"),
   647 => (x"72",x"87",x"c2",x"79"),
   648 => (x"02",x"9c",x"74",x"8c"),
   649 => (x"1e",x"49",x"87",x"dd"),
   650 => (x"fb",x"fa",x"49",x"73"),
   651 => (x"d4",x"86",x"c4",x"87"),
   652 => (x"ff",x"c7",x"49",x"66"),
   653 => (x"87",x"cb",x"02",x"99"),
   654 => (x"1e",x"de",x"f5",x"c2"),
   655 => (x"c1",x"fc",x"49",x"73"),
   656 => (x"26",x"86",x"c4",x"87"),
   657 => (x"1e",x"87",x"cd",x"f5"),
   658 => (x"4b",x"71",x"1e",x"73"),
   659 => (x"e4",x"c0",x"02",x"9b"),
   660 => (x"cb",x"c2",x"c3",x"87"),
   661 => (x"c2",x"4a",x"73",x"5b"),
   662 => (x"de",x"fd",x"c2",x"8a"),
   663 => (x"c3",x"92",x"49",x"bf"),
   664 => (x"48",x"bf",x"f7",x"c1"),
   665 => (x"c2",x"c3",x"80",x"72"),
   666 => (x"48",x"71",x"58",x"cf"),
   667 => (x"fd",x"c2",x"30",x"c4"),
   668 => (x"ed",x"c0",x"58",x"ee"),
   669 => (x"c7",x"c2",x"c3",x"87"),
   670 => (x"fb",x"c1",x"c3",x"48"),
   671 => (x"c2",x"c3",x"78",x"bf"),
   672 => (x"c1",x"c3",x"48",x"cb"),
   673 => (x"c2",x"78",x"bf",x"ff"),
   674 => (x"02",x"bf",x"e6",x"fd"),
   675 => (x"fd",x"c2",x"87",x"c9"),
   676 => (x"c4",x"49",x"bf",x"de"),
   677 => (x"c3",x"87",x"c7",x"31"),
   678 => (x"49",x"bf",x"c3",x"c2"),
   679 => (x"fd",x"c2",x"31",x"c4"),
   680 => (x"f3",x"f3",x"59",x"ee"),
   681 => (x"5b",x"5e",x"0e",x"87"),
   682 => (x"4a",x"71",x"0e",x"5c"),
   683 => (x"9a",x"72",x"4b",x"c0"),
   684 => (x"87",x"e1",x"c0",x"02"),
   685 => (x"9f",x"49",x"a2",x"da"),
   686 => (x"fd",x"c2",x"4b",x"69"),
   687 => (x"cf",x"02",x"bf",x"e6"),
   688 => (x"49",x"a2",x"d4",x"87"),
   689 => (x"4c",x"49",x"69",x"9f"),
   690 => (x"9c",x"ff",x"ff",x"c0"),
   691 => (x"87",x"c2",x"34",x"d0"),
   692 => (x"49",x"74",x"4c",x"c0"),
   693 => (x"fd",x"49",x"73",x"b3"),
   694 => (x"f9",x"f2",x"87",x"ed"),
   695 => (x"5b",x"5e",x"0e",x"87"),
   696 => (x"f4",x"0e",x"5d",x"5c"),
   697 => (x"c0",x"4a",x"71",x"86"),
   698 => (x"02",x"9a",x"72",x"7e"),
   699 => (x"f5",x"c2",x"87",x"d8"),
   700 => (x"78",x"c0",x"48",x"da"),
   701 => (x"48",x"d2",x"f5",x"c2"),
   702 => (x"bf",x"cb",x"c2",x"c3"),
   703 => (x"d6",x"f5",x"c2",x"78"),
   704 => (x"c7",x"c2",x"c3",x"48"),
   705 => (x"fd",x"c2",x"78",x"bf"),
   706 => (x"50",x"c0",x"48",x"fb"),
   707 => (x"bf",x"ea",x"fd",x"c2"),
   708 => (x"da",x"f5",x"c2",x"49"),
   709 => (x"aa",x"71",x"4a",x"bf"),
   710 => (x"87",x"c9",x"c4",x"03"),
   711 => (x"99",x"cf",x"49",x"72"),
   712 => (x"87",x"e9",x"c0",x"05"),
   713 => (x"48",x"f8",x"f2",x"c0"),
   714 => (x"bf",x"d2",x"f5",x"c2"),
   715 => (x"de",x"f5",x"c2",x"78"),
   716 => (x"d2",x"f5",x"c2",x"1e"),
   717 => (x"f5",x"c2",x"49",x"bf"),
   718 => (x"a1",x"c1",x"48",x"d2"),
   719 => (x"d5",x"e3",x"71",x"78"),
   720 => (x"c0",x"86",x"c4",x"87"),
   721 => (x"c2",x"48",x"f4",x"f2"),
   722 => (x"cc",x"78",x"de",x"f5"),
   723 => (x"f4",x"f2",x"c0",x"87"),
   724 => (x"e0",x"c0",x"48",x"bf"),
   725 => (x"f8",x"f2",x"c0",x"80"),
   726 => (x"da",x"f5",x"c2",x"58"),
   727 => (x"80",x"c1",x"48",x"bf"),
   728 => (x"58",x"de",x"f5",x"c2"),
   729 => (x"00",x"0c",x"b4",x"27"),
   730 => (x"bf",x"97",x"bf",x"00"),
   731 => (x"c2",x"02",x"9d",x"4d"),
   732 => (x"e5",x"c3",x"87",x"e3"),
   733 => (x"dc",x"c2",x"02",x"ad"),
   734 => (x"f4",x"f2",x"c0",x"87"),
   735 => (x"a3",x"cb",x"4b",x"bf"),
   736 => (x"cf",x"4c",x"11",x"49"),
   737 => (x"d2",x"c1",x"05",x"ac"),
   738 => (x"df",x"49",x"75",x"87"),
   739 => (x"cd",x"89",x"c1",x"99"),
   740 => (x"ee",x"fd",x"c2",x"91"),
   741 => (x"4a",x"a3",x"c1",x"81"),
   742 => (x"a3",x"c3",x"51",x"12"),
   743 => (x"c5",x"51",x"12",x"4a"),
   744 => (x"51",x"12",x"4a",x"a3"),
   745 => (x"12",x"4a",x"a3",x"c7"),
   746 => (x"4a",x"a3",x"c9",x"51"),
   747 => (x"a3",x"ce",x"51",x"12"),
   748 => (x"d0",x"51",x"12",x"4a"),
   749 => (x"51",x"12",x"4a",x"a3"),
   750 => (x"12",x"4a",x"a3",x"d2"),
   751 => (x"4a",x"a3",x"d4",x"51"),
   752 => (x"a3",x"d6",x"51",x"12"),
   753 => (x"d8",x"51",x"12",x"4a"),
   754 => (x"51",x"12",x"4a",x"a3"),
   755 => (x"12",x"4a",x"a3",x"dc"),
   756 => (x"4a",x"a3",x"de",x"51"),
   757 => (x"7e",x"c1",x"51",x"12"),
   758 => (x"74",x"87",x"fa",x"c0"),
   759 => (x"05",x"99",x"c8",x"49"),
   760 => (x"74",x"87",x"eb",x"c0"),
   761 => (x"05",x"99",x"d0",x"49"),
   762 => (x"66",x"dc",x"87",x"d1"),
   763 => (x"87",x"cb",x"c0",x"02"),
   764 => (x"66",x"dc",x"49",x"73"),
   765 => (x"02",x"98",x"70",x"0f"),
   766 => (x"6e",x"87",x"d3",x"c0"),
   767 => (x"87",x"c6",x"c0",x"05"),
   768 => (x"48",x"ee",x"fd",x"c2"),
   769 => (x"f2",x"c0",x"50",x"c0"),
   770 => (x"c2",x"48",x"bf",x"f4"),
   771 => (x"fd",x"c2",x"87",x"e1"),
   772 => (x"50",x"c0",x"48",x"fb"),
   773 => (x"ea",x"fd",x"c2",x"7e"),
   774 => (x"f5",x"c2",x"49",x"bf"),
   775 => (x"71",x"4a",x"bf",x"da"),
   776 => (x"f7",x"fb",x"04",x"aa"),
   777 => (x"cb",x"c2",x"c3",x"87"),
   778 => (x"c8",x"c0",x"05",x"bf"),
   779 => (x"e6",x"fd",x"c2",x"87"),
   780 => (x"f8",x"c1",x"02",x"bf"),
   781 => (x"d6",x"f5",x"c2",x"87"),
   782 => (x"df",x"ed",x"49",x"bf"),
   783 => (x"c2",x"49",x"70",x"87"),
   784 => (x"c4",x"59",x"da",x"f5"),
   785 => (x"f5",x"c2",x"48",x"a6"),
   786 => (x"c2",x"78",x"bf",x"d6"),
   787 => (x"02",x"bf",x"e6",x"fd"),
   788 => (x"c4",x"87",x"d8",x"c0"),
   789 => (x"ff",x"cf",x"49",x"66"),
   790 => (x"99",x"f8",x"ff",x"ff"),
   791 => (x"c5",x"c0",x"02",x"a9"),
   792 => (x"c0",x"4c",x"c0",x"87"),
   793 => (x"4c",x"c1",x"87",x"e1"),
   794 => (x"c4",x"87",x"dc",x"c0"),
   795 => (x"ff",x"cf",x"49",x"66"),
   796 => (x"02",x"a9",x"99",x"f8"),
   797 => (x"c8",x"87",x"c8",x"c0"),
   798 => (x"78",x"c0",x"48",x"a6"),
   799 => (x"c8",x"87",x"c5",x"c0"),
   800 => (x"78",x"c1",x"48",x"a6"),
   801 => (x"74",x"4c",x"66",x"c8"),
   802 => (x"e0",x"c0",x"05",x"9c"),
   803 => (x"49",x"66",x"c4",x"87"),
   804 => (x"fd",x"c2",x"89",x"c2"),
   805 => (x"91",x"4a",x"bf",x"de"),
   806 => (x"bf",x"f7",x"c1",x"c3"),
   807 => (x"d2",x"f5",x"c2",x"4a"),
   808 => (x"78",x"a1",x"72",x"48"),
   809 => (x"48",x"da",x"f5",x"c2"),
   810 => (x"df",x"f9",x"78",x"c0"),
   811 => (x"f4",x"48",x"c0",x"87"),
   812 => (x"87",x"e0",x"eb",x"8e"),
   813 => (x"00",x"00",x"00",x"00"),
   814 => (x"ff",x"ff",x"ff",x"ff"),
   815 => (x"00",x"00",x"0c",x"c4"),
   816 => (x"00",x"00",x"0c",x"cd"),
   817 => (x"33",x"54",x"41",x"46"),
   818 => (x"20",x"20",x"20",x"32"),
   819 => (x"54",x"41",x"46",x"00"),
   820 => (x"20",x"20",x"36",x"31"),
   821 => (x"ff",x"1e",x"00",x"20"),
   822 => (x"ff",x"c3",x"48",x"d4"),
   823 => (x"26",x"48",x"68",x"78"),
   824 => (x"d4",x"ff",x"1e",x"4f"),
   825 => (x"78",x"ff",x"c3",x"48"),
   826 => (x"c8",x"48",x"d0",x"ff"),
   827 => (x"d4",x"ff",x"78",x"e1"),
   828 => (x"c3",x"78",x"d4",x"48"),
   829 => (x"ff",x"48",x"cf",x"c2"),
   830 => (x"26",x"50",x"bf",x"d4"),
   831 => (x"d0",x"ff",x"1e",x"4f"),
   832 => (x"78",x"e0",x"c0",x"48"),
   833 => (x"ff",x"1e",x"4f",x"26"),
   834 => (x"49",x"70",x"87",x"cc"),
   835 => (x"87",x"c6",x"02",x"99"),
   836 => (x"05",x"a9",x"fb",x"c0"),
   837 => (x"48",x"71",x"87",x"f1"),
   838 => (x"5e",x"0e",x"4f",x"26"),
   839 => (x"71",x"0e",x"5c",x"5b"),
   840 => (x"fe",x"4c",x"c0",x"4b"),
   841 => (x"49",x"70",x"87",x"f0"),
   842 => (x"f9",x"c0",x"02",x"99"),
   843 => (x"a9",x"ec",x"c0",x"87"),
   844 => (x"87",x"f2",x"c0",x"02"),
   845 => (x"02",x"a9",x"fb",x"c0"),
   846 => (x"cc",x"87",x"eb",x"c0"),
   847 => (x"03",x"ac",x"b7",x"66"),
   848 => (x"66",x"d0",x"87",x"c7"),
   849 => (x"71",x"87",x"c2",x"02"),
   850 => (x"02",x"99",x"71",x"53"),
   851 => (x"84",x"c1",x"87",x"c2"),
   852 => (x"70",x"87",x"c3",x"fe"),
   853 => (x"cd",x"02",x"99",x"49"),
   854 => (x"a9",x"ec",x"c0",x"87"),
   855 => (x"c0",x"87",x"c7",x"02"),
   856 => (x"ff",x"05",x"a9",x"fb"),
   857 => (x"66",x"d0",x"87",x"d5"),
   858 => (x"c0",x"87",x"c3",x"02"),
   859 => (x"ec",x"c0",x"7b",x"97"),
   860 => (x"87",x"c4",x"05",x"a9"),
   861 => (x"87",x"c5",x"4a",x"74"),
   862 => (x"0a",x"c0",x"4a",x"74"),
   863 => (x"c2",x"48",x"72",x"8a"),
   864 => (x"26",x"4d",x"26",x"87"),
   865 => (x"26",x"4b",x"26",x"4c"),
   866 => (x"c9",x"fd",x"1e",x"4f"),
   867 => (x"c0",x"49",x"70",x"87"),
   868 => (x"04",x"a9",x"b7",x"f0"),
   869 => (x"f9",x"c0",x"87",x"ca"),
   870 => (x"c3",x"01",x"a9",x"b7"),
   871 => (x"89",x"f0",x"c0",x"87"),
   872 => (x"a9",x"b7",x"c1",x"c1"),
   873 => (x"c1",x"87",x"ca",x"04"),
   874 => (x"01",x"a9",x"b7",x"da"),
   875 => (x"f7",x"c0",x"87",x"c3"),
   876 => (x"b7",x"e1",x"c1",x"89"),
   877 => (x"87",x"ca",x"04",x"a9"),
   878 => (x"a9",x"b7",x"fa",x"c1"),
   879 => (x"c0",x"87",x"c3",x"01"),
   880 => (x"48",x"71",x"89",x"fd"),
   881 => (x"5e",x"0e",x"4f",x"26"),
   882 => (x"71",x"0e",x"5c",x"5b"),
   883 => (x"4c",x"d4",x"ff",x"4a"),
   884 => (x"ea",x"c0",x"49",x"72"),
   885 => (x"9b",x"4b",x"70",x"87"),
   886 => (x"c1",x"87",x"c2",x"02"),
   887 => (x"48",x"d0",x"ff",x"8b"),
   888 => (x"c1",x"78",x"c5",x"c8"),
   889 => (x"49",x"73",x"7c",x"d5"),
   890 => (x"e7",x"c1",x"31",x"c6"),
   891 => (x"4a",x"bf",x"97",x"e5"),
   892 => (x"70",x"b0",x"71",x"48"),
   893 => (x"48",x"d0",x"ff",x"7c"),
   894 => (x"48",x"73",x"78",x"c4"),
   895 => (x"0e",x"87",x"c4",x"fe"),
   896 => (x"5d",x"5c",x"5b",x"5e"),
   897 => (x"71",x"86",x"f8",x"0e"),
   898 => (x"c0",x"7e",x"c0",x"4b"),
   899 => (x"bf",x"97",x"e6",x"fb"),
   900 => (x"05",x"a9",x"df",x"49"),
   901 => (x"c8",x"87",x"ee",x"c0"),
   902 => (x"69",x"97",x"49",x"a3"),
   903 => (x"a9",x"c3",x"c1",x"49"),
   904 => (x"c9",x"87",x"dd",x"05"),
   905 => (x"69",x"97",x"49",x"a3"),
   906 => (x"a9",x"c6",x"c1",x"49"),
   907 => (x"ca",x"87",x"d1",x"05"),
   908 => (x"69",x"97",x"49",x"a3"),
   909 => (x"a9",x"c7",x"c1",x"49"),
   910 => (x"c1",x"87",x"c5",x"05"),
   911 => (x"87",x"e1",x"c2",x"48"),
   912 => (x"dc",x"c2",x"48",x"c0"),
   913 => (x"87",x"d9",x"fa",x"87"),
   914 => (x"fb",x"c0",x"4c",x"c0"),
   915 => (x"49",x"bf",x"97",x"e6"),
   916 => (x"cf",x"04",x"a9",x"c0"),
   917 => (x"87",x"ee",x"fa",x"87"),
   918 => (x"fb",x"c0",x"84",x"c1"),
   919 => (x"49",x"bf",x"97",x"e6"),
   920 => (x"87",x"f1",x"06",x"ac"),
   921 => (x"97",x"e6",x"fb",x"c0"),
   922 => (x"87",x"cf",x"02",x"bf"),
   923 => (x"70",x"87",x"e7",x"f9"),
   924 => (x"c6",x"02",x"99",x"49"),
   925 => (x"a9",x"ec",x"c0",x"87"),
   926 => (x"c0",x"87",x"f1",x"05"),
   927 => (x"87",x"d6",x"f9",x"4c"),
   928 => (x"d1",x"f9",x"4d",x"70"),
   929 => (x"58",x"a6",x"c8",x"87"),
   930 => (x"70",x"87",x"cb",x"f9"),
   931 => (x"c8",x"84",x"c1",x"4a"),
   932 => (x"69",x"97",x"49",x"a3"),
   933 => (x"c7",x"02",x"ad",x"49"),
   934 => (x"ad",x"ff",x"c0",x"87"),
   935 => (x"87",x"e7",x"c0",x"05"),
   936 => (x"97",x"49",x"a3",x"c9"),
   937 => (x"66",x"c4",x"49",x"69"),
   938 => (x"87",x"c7",x"02",x"a9"),
   939 => (x"a8",x"ff",x"c0",x"48"),
   940 => (x"ca",x"87",x"d4",x"05"),
   941 => (x"69",x"97",x"49",x"a3"),
   942 => (x"c6",x"02",x"aa",x"49"),
   943 => (x"aa",x"ff",x"c0",x"87"),
   944 => (x"c1",x"87",x"c4",x"05"),
   945 => (x"c0",x"87",x"d0",x"7e"),
   946 => (x"c6",x"02",x"ad",x"ec"),
   947 => (x"ad",x"fb",x"c0",x"87"),
   948 => (x"c0",x"87",x"c4",x"05"),
   949 => (x"6e",x"7e",x"c1",x"4c"),
   950 => (x"87",x"e1",x"fe",x"02"),
   951 => (x"74",x"87",x"de",x"f8"),
   952 => (x"fa",x"8e",x"f8",x"48"),
   953 => (x"0e",x"00",x"87",x"db"),
   954 => (x"5d",x"5c",x"5b",x"5e"),
   955 => (x"4d",x"71",x"1e",x"0e"),
   956 => (x"75",x"4b",x"d4",x"ff"),
   957 => (x"d4",x"c2",x"c3",x"1e"),
   958 => (x"87",x"f1",x"e5",x"49"),
   959 => (x"98",x"70",x"86",x"c4"),
   960 => (x"87",x"d8",x"c3",x"02"),
   961 => (x"bf",x"dc",x"c2",x"c3"),
   962 => (x"fa",x"49",x"75",x"4c"),
   963 => (x"d0",x"ff",x"87",x"f8"),
   964 => (x"78",x"c5",x"c8",x"48"),
   965 => (x"c0",x"7b",x"d6",x"c1"),
   966 => (x"49",x"a2",x"75",x"4a"),
   967 => (x"82",x"c1",x"7b",x"11"),
   968 => (x"04",x"aa",x"b7",x"cb"),
   969 => (x"4a",x"cc",x"87",x"f3"),
   970 => (x"c1",x"7b",x"ff",x"c3"),
   971 => (x"b7",x"e0",x"c0",x"82"),
   972 => (x"87",x"f4",x"04",x"aa"),
   973 => (x"c4",x"48",x"d0",x"ff"),
   974 => (x"7b",x"ff",x"c3",x"78"),
   975 => (x"c1",x"78",x"c5",x"c8"),
   976 => (x"7b",x"c1",x"7b",x"d3"),
   977 => (x"9c",x"74",x"78",x"c4"),
   978 => (x"87",x"ff",x"c1",x"02"),
   979 => (x"7e",x"de",x"f5",x"c2"),
   980 => (x"8c",x"4d",x"c0",x"c8"),
   981 => (x"03",x"ac",x"b7",x"c0"),
   982 => (x"c0",x"c8",x"87",x"c6"),
   983 => (x"4c",x"c0",x"4d",x"a4"),
   984 => (x"05",x"ad",x"c0",x"c8"),
   985 => (x"c2",x"c3",x"87",x"dc"),
   986 => (x"49",x"bf",x"97",x"cf"),
   987 => (x"d1",x"02",x"99",x"d0"),
   988 => (x"c3",x"1e",x"c0",x"87"),
   989 => (x"e7",x"49",x"d4",x"c2"),
   990 => (x"86",x"c4",x"87",x"c8"),
   991 => (x"c0",x"4a",x"49",x"70"),
   992 => (x"f5",x"c2",x"87",x"ee"),
   993 => (x"c2",x"c3",x"1e",x"de"),
   994 => (x"f5",x"e6",x"49",x"d4"),
   995 => (x"70",x"86",x"c4",x"87"),
   996 => (x"d0",x"ff",x"4a",x"49"),
   997 => (x"78",x"c5",x"c8",x"48"),
   998 => (x"6e",x"7b",x"d4",x"c1"),
   999 => (x"6e",x"7b",x"bf",x"97"),
  1000 => (x"70",x"80",x"c1",x"48"),
  1001 => (x"05",x"8d",x"c1",x"7e"),
  1002 => (x"ff",x"87",x"f0",x"ff"),
  1003 => (x"78",x"c4",x"48",x"d0"),
  1004 => (x"c5",x"05",x"9a",x"72"),
  1005 => (x"c0",x"48",x"c0",x"87"),
  1006 => (x"1e",x"c1",x"87",x"e4"),
  1007 => (x"49",x"d4",x"c2",x"c3"),
  1008 => (x"c4",x"87",x"e5",x"e4"),
  1009 => (x"05",x"9c",x"74",x"86"),
  1010 => (x"ff",x"87",x"c1",x"fe"),
  1011 => (x"c5",x"c8",x"48",x"d0"),
  1012 => (x"7b",x"d3",x"c1",x"78"),
  1013 => (x"78",x"c4",x"7b",x"c0"),
  1014 => (x"87",x"c2",x"48",x"c1"),
  1015 => (x"26",x"26",x"48",x"c0"),
  1016 => (x"26",x"4c",x"26",x"4d"),
  1017 => (x"0e",x"4f",x"26",x"4b"),
  1018 => (x"5d",x"5c",x"5b",x"5e"),
  1019 => (x"4b",x"71",x"1e",x"0e"),
  1020 => (x"ab",x"4d",x"4c",x"c0"),
  1021 => (x"87",x"e8",x"c0",x"04"),
  1022 => (x"1e",x"ff",x"f7",x"c0"),
  1023 => (x"c4",x"02",x"9d",x"75"),
  1024 => (x"c2",x"4a",x"c0",x"87"),
  1025 => (x"72",x"4a",x"c1",x"87"),
  1026 => (x"87",x"d1",x"eb",x"49"),
  1027 => (x"7e",x"70",x"86",x"c4"),
  1028 => (x"05",x"6e",x"84",x"c1"),
  1029 => (x"4c",x"73",x"87",x"c2"),
  1030 => (x"ac",x"73",x"85",x"c1"),
  1031 => (x"87",x"d8",x"ff",x"06"),
  1032 => (x"fe",x"26",x"48",x"6e"),
  1033 => (x"5e",x"0e",x"87",x"f9"),
  1034 => (x"71",x"0e",x"5c",x"5b"),
  1035 => (x"02",x"66",x"cc",x"4b"),
  1036 => (x"4c",x"87",x"e8",x"c0"),
  1037 => (x"02",x"8c",x"f0",x"c0"),
  1038 => (x"74",x"87",x"e8",x"c0"),
  1039 => (x"02",x"8a",x"c1",x"4a"),
  1040 => (x"8a",x"87",x"e0",x"c0"),
  1041 => (x"8a",x"87",x"dc",x"02"),
  1042 => (x"c0",x"87",x"d8",x"02"),
  1043 => (x"c0",x"02",x"8a",x"e0"),
  1044 => (x"8a",x"c1",x"87",x"e5"),
  1045 => (x"87",x"e7",x"c0",x"02"),
  1046 => (x"73",x"87",x"ea",x"c0"),
  1047 => (x"87",x"c7",x"fa",x"49"),
  1048 => (x"74",x"87",x"e2",x"c0"),
  1049 => (x"c1",x"49",x"c0",x"1e"),
  1050 => (x"74",x"87",x"d7",x"ed"),
  1051 => (x"c1",x"49",x"73",x"1e"),
  1052 => (x"c8",x"87",x"cf",x"ed"),
  1053 => (x"73",x"87",x"ce",x"86"),
  1054 => (x"c5",x"f1",x"c1",x"49"),
  1055 => (x"73",x"87",x"c6",x"87"),
  1056 => (x"f5",x"f1",x"c1",x"49"),
  1057 => (x"87",x"d9",x"fd",x"87"),
  1058 => (x"5c",x"5b",x"5e",x"0e"),
  1059 => (x"71",x"1e",x"0e",x"5d"),
  1060 => (x"91",x"de",x"49",x"4c"),
  1061 => (x"4d",x"fc",x"c2",x"c3"),
  1062 => (x"6d",x"97",x"85",x"71"),
  1063 => (x"87",x"dc",x"c1",x"02"),
  1064 => (x"bf",x"e8",x"c2",x"c3"),
  1065 => (x"72",x"82",x"74",x"4a"),
  1066 => (x"87",x"fb",x"fc",x"49"),
  1067 => (x"02",x"6e",x"7e",x"70"),
  1068 => (x"c3",x"87",x"f2",x"c0"),
  1069 => (x"6e",x"4b",x"f0",x"c2"),
  1070 => (x"fe",x"49",x"cb",x"4a"),
  1071 => (x"74",x"87",x"e9",x"ff"),
  1072 => (x"c1",x"93",x"cb",x"4b"),
  1073 => (x"c4",x"83",x"d8",x"e8"),
  1074 => (x"c0",x"c4",x"c1",x"83"),
  1075 => (x"c1",x"49",x"74",x"7b"),
  1076 => (x"75",x"87",x"fa",x"d6"),
  1077 => (x"e6",x"e7",x"c1",x"7b"),
  1078 => (x"1e",x"49",x"bf",x"97"),
  1079 => (x"49",x"f0",x"c2",x"c3"),
  1080 => (x"c4",x"87",x"c3",x"fd"),
  1081 => (x"c1",x"49",x"74",x"86"),
  1082 => (x"c0",x"87",x"e2",x"d6"),
  1083 => (x"c1",x"d8",x"c1",x"49"),
  1084 => (x"d0",x"c2",x"c3",x"87"),
  1085 => (x"c1",x"78",x"c0",x"48"),
  1086 => (x"87",x"f0",x"df",x"49"),
  1087 => (x"87",x"df",x"fb",x"26"),
  1088 => (x"64",x"61",x"6f",x"4c"),
  1089 => (x"2e",x"67",x"6e",x"69"),
  1090 => (x"0e",x"00",x"2e",x"2e"),
  1091 => (x"0e",x"5c",x"5b",x"5e"),
  1092 => (x"c3",x"4a",x"4b",x"71"),
  1093 => (x"82",x"bf",x"e8",x"c2"),
  1094 => (x"ca",x"fb",x"49",x"72"),
  1095 => (x"9c",x"4c",x"70",x"87"),
  1096 => (x"49",x"87",x"c4",x"02"),
  1097 => (x"c3",x"87",x"fe",x"e5"),
  1098 => (x"c0",x"48",x"e8",x"c2"),
  1099 => (x"de",x"49",x"c1",x"78"),
  1100 => (x"ec",x"fa",x"87",x"fa"),
  1101 => (x"5b",x"5e",x"0e",x"87"),
  1102 => (x"f4",x"0e",x"5d",x"5c"),
  1103 => (x"de",x"f5",x"c2",x"86"),
  1104 => (x"c4",x"4c",x"c0",x"4d"),
  1105 => (x"78",x"c0",x"48",x"a6"),
  1106 => (x"bf",x"e8",x"c2",x"c3"),
  1107 => (x"06",x"a9",x"c0",x"49"),
  1108 => (x"c2",x"87",x"c1",x"c1"),
  1109 => (x"98",x"48",x"de",x"f5"),
  1110 => (x"87",x"f8",x"c0",x"02"),
  1111 => (x"1e",x"ff",x"f7",x"c0"),
  1112 => (x"c7",x"02",x"66",x"c8"),
  1113 => (x"48",x"a6",x"c4",x"87"),
  1114 => (x"87",x"c5",x"78",x"c0"),
  1115 => (x"c1",x"48",x"a6",x"c4"),
  1116 => (x"49",x"66",x"c4",x"78"),
  1117 => (x"c4",x"87",x"e6",x"e5"),
  1118 => (x"c1",x"4d",x"70",x"86"),
  1119 => (x"48",x"66",x"c4",x"84"),
  1120 => (x"a6",x"c8",x"80",x"c1"),
  1121 => (x"e8",x"c2",x"c3",x"58"),
  1122 => (x"03",x"ac",x"49",x"bf"),
  1123 => (x"9d",x"75",x"87",x"c6"),
  1124 => (x"87",x"c8",x"ff",x"05"),
  1125 => (x"9d",x"75",x"4c",x"c0"),
  1126 => (x"87",x"e0",x"c3",x"02"),
  1127 => (x"1e",x"ff",x"f7",x"c0"),
  1128 => (x"c7",x"02",x"66",x"c8"),
  1129 => (x"48",x"a6",x"cc",x"87"),
  1130 => (x"87",x"c5",x"78",x"c0"),
  1131 => (x"c1",x"48",x"a6",x"cc"),
  1132 => (x"49",x"66",x"cc",x"78"),
  1133 => (x"c4",x"87",x"e6",x"e4"),
  1134 => (x"6e",x"7e",x"70",x"86"),
  1135 => (x"87",x"e9",x"c2",x"02"),
  1136 => (x"81",x"cb",x"49",x"6e"),
  1137 => (x"d0",x"49",x"69",x"97"),
  1138 => (x"d6",x"c1",x"02",x"99"),
  1139 => (x"cb",x"c4",x"c1",x"87"),
  1140 => (x"cb",x"49",x"74",x"4a"),
  1141 => (x"d8",x"e8",x"c1",x"91"),
  1142 => (x"c8",x"79",x"72",x"81"),
  1143 => (x"51",x"ff",x"c3",x"81"),
  1144 => (x"91",x"de",x"49",x"74"),
  1145 => (x"4d",x"fc",x"c2",x"c3"),
  1146 => (x"c1",x"c2",x"85",x"71"),
  1147 => (x"a5",x"c1",x"7d",x"97"),
  1148 => (x"51",x"e0",x"c0",x"49"),
  1149 => (x"97",x"ee",x"fd",x"c2"),
  1150 => (x"87",x"d2",x"02",x"bf"),
  1151 => (x"a5",x"c2",x"84",x"c1"),
  1152 => (x"ee",x"fd",x"c2",x"4b"),
  1153 => (x"fe",x"49",x"db",x"4a"),
  1154 => (x"c1",x"87",x"dd",x"fa"),
  1155 => (x"a5",x"cd",x"87",x"db"),
  1156 => (x"c1",x"51",x"c0",x"49"),
  1157 => (x"4b",x"a5",x"c2",x"84"),
  1158 => (x"49",x"cb",x"4a",x"6e"),
  1159 => (x"87",x"c8",x"fa",x"fe"),
  1160 => (x"c1",x"87",x"c6",x"c1"),
  1161 => (x"74",x"4a",x"c8",x"c2"),
  1162 => (x"c1",x"91",x"cb",x"49"),
  1163 => (x"72",x"81",x"d8",x"e8"),
  1164 => (x"ee",x"fd",x"c2",x"79"),
  1165 => (x"d8",x"02",x"bf",x"97"),
  1166 => (x"de",x"49",x"74",x"87"),
  1167 => (x"c3",x"84",x"c1",x"91"),
  1168 => (x"71",x"4b",x"fc",x"c2"),
  1169 => (x"ee",x"fd",x"c2",x"83"),
  1170 => (x"fe",x"49",x"dd",x"4a"),
  1171 => (x"d8",x"87",x"d9",x"f9"),
  1172 => (x"de",x"4b",x"74",x"87"),
  1173 => (x"fc",x"c2",x"c3",x"93"),
  1174 => (x"49",x"a3",x"cb",x"83"),
  1175 => (x"84",x"c1",x"51",x"c0"),
  1176 => (x"cb",x"4a",x"6e",x"73"),
  1177 => (x"ff",x"f8",x"fe",x"49"),
  1178 => (x"48",x"66",x"c4",x"87"),
  1179 => (x"a6",x"c8",x"80",x"c1"),
  1180 => (x"03",x"ac",x"c7",x"58"),
  1181 => (x"6e",x"87",x"c5",x"c0"),
  1182 => (x"87",x"e0",x"fc",x"05"),
  1183 => (x"8e",x"f4",x"48",x"74"),
  1184 => (x"1e",x"87",x"dc",x"f5"),
  1185 => (x"4b",x"71",x"1e",x"73"),
  1186 => (x"c1",x"91",x"cb",x"49"),
  1187 => (x"c8",x"81",x"d8",x"e8"),
  1188 => (x"e7",x"c1",x"4a",x"a1"),
  1189 => (x"50",x"12",x"48",x"e5"),
  1190 => (x"c0",x"4a",x"a1",x"c9"),
  1191 => (x"12",x"48",x"e6",x"fb"),
  1192 => (x"c1",x"81",x"ca",x"50"),
  1193 => (x"11",x"48",x"e6",x"e7"),
  1194 => (x"e6",x"e7",x"c1",x"50"),
  1195 => (x"1e",x"49",x"bf",x"97"),
  1196 => (x"f1",x"f5",x"49",x"c0"),
  1197 => (x"d0",x"c2",x"c3",x"87"),
  1198 => (x"c1",x"78",x"de",x"48"),
  1199 => (x"87",x"ec",x"d8",x"49"),
  1200 => (x"87",x"df",x"f4",x"26"),
  1201 => (x"49",x"4a",x"71",x"1e"),
  1202 => (x"e8",x"c1",x"91",x"cb"),
  1203 => (x"81",x"c8",x"81",x"d8"),
  1204 => (x"c2",x"c3",x"48",x"11"),
  1205 => (x"c2",x"c3",x"58",x"d4"),
  1206 => (x"78",x"c0",x"48",x"e8"),
  1207 => (x"cb",x"d8",x"49",x"c1"),
  1208 => (x"1e",x"4f",x"26",x"87"),
  1209 => (x"d0",x"c1",x"49",x"c0"),
  1210 => (x"4f",x"26",x"87",x"c8"),
  1211 => (x"02",x"99",x"71",x"1e"),
  1212 => (x"e9",x"c1",x"87",x"d2"),
  1213 => (x"50",x"c0",x"48",x"ed"),
  1214 => (x"cb",x"c1",x"80",x"f7"),
  1215 => (x"e8",x"c1",x"40",x"c4"),
  1216 => (x"87",x"ce",x"78",x"c6"),
  1217 => (x"48",x"e9",x"e9",x"c1"),
  1218 => (x"78",x"e7",x"e7",x"c1"),
  1219 => (x"cb",x"c1",x"80",x"fc"),
  1220 => (x"4f",x"26",x"78",x"e3"),
  1221 => (x"5c",x"5b",x"5e",x"0e"),
  1222 => (x"4a",x"4c",x"71",x"0e"),
  1223 => (x"e8",x"c1",x"92",x"cb"),
  1224 => (x"a2",x"c8",x"82",x"d8"),
  1225 => (x"4b",x"a2",x"c9",x"49"),
  1226 => (x"1e",x"4b",x"6b",x"97"),
  1227 => (x"1e",x"49",x"69",x"97"),
  1228 => (x"49",x"12",x"82",x"ca"),
  1229 => (x"87",x"c1",x"f9",x"c0"),
  1230 => (x"ef",x"d6",x"49",x"c0"),
  1231 => (x"c1",x"49",x"74",x"87"),
  1232 => (x"f8",x"87",x"ca",x"cd"),
  1233 => (x"87",x"d9",x"f2",x"8e"),
  1234 => (x"71",x"1e",x"73",x"1e"),
  1235 => (x"c3",x"ff",x"49",x"4b"),
  1236 => (x"fe",x"49",x"73",x"87"),
  1237 => (x"ca",x"f2",x"87",x"fe"),
  1238 => (x"1e",x"73",x"1e",x"87"),
  1239 => (x"a3",x"c6",x"4b",x"71"),
  1240 => (x"87",x"dc",x"02",x"4a"),
  1241 => (x"c0",x"02",x"8a",x"c1"),
  1242 => (x"02",x"8a",x"87",x"e4"),
  1243 => (x"8a",x"87",x"e8",x"c1"),
  1244 => (x"87",x"ca",x"c1",x"02"),
  1245 => (x"ef",x"c0",x"02",x"8a"),
  1246 => (x"d9",x"02",x"8a",x"87"),
  1247 => (x"87",x"e9",x"c1",x"87"),
  1248 => (x"48",x"d0",x"c2",x"c3"),
  1249 => (x"49",x"c1",x"78",x"df"),
  1250 => (x"c1",x"87",x"e1",x"d5"),
  1251 => (x"49",x"c7",x"87",x"e6"),
  1252 => (x"c1",x"87",x"f1",x"fc"),
  1253 => (x"c2",x"c3",x"87",x"de"),
  1254 => (x"c1",x"02",x"bf",x"e8"),
  1255 => (x"c1",x"48",x"87",x"cb"),
  1256 => (x"ec",x"c2",x"c3",x"88"),
  1257 => (x"87",x"c1",x"c1",x"58"),
  1258 => (x"bf",x"ec",x"c2",x"c3"),
  1259 => (x"87",x"f9",x"c0",x"02"),
  1260 => (x"bf",x"e8",x"c2",x"c3"),
  1261 => (x"c3",x"80",x"c1",x"48"),
  1262 => (x"c0",x"58",x"ec",x"c2"),
  1263 => (x"c2",x"c3",x"87",x"eb"),
  1264 => (x"c6",x"49",x"bf",x"e8"),
  1265 => (x"ec",x"c2",x"c3",x"89"),
  1266 => (x"a9",x"b7",x"c0",x"59"),
  1267 => (x"c3",x"87",x"da",x"03"),
  1268 => (x"c0",x"48",x"e8",x"c2"),
  1269 => (x"c3",x"87",x"d2",x"78"),
  1270 => (x"02",x"bf",x"ec",x"c2"),
  1271 => (x"c2",x"c3",x"87",x"cb"),
  1272 => (x"c6",x"48",x"bf",x"e8"),
  1273 => (x"ec",x"c2",x"c3",x"80"),
  1274 => (x"d3",x"49",x"c0",x"58"),
  1275 => (x"49",x"73",x"87",x"fe"),
  1276 => (x"87",x"d9",x"ca",x"c1"),
  1277 => (x"0e",x"87",x"ec",x"ef"),
  1278 => (x"0e",x"5c",x"5b",x"5e"),
  1279 => (x"66",x"cc",x"4c",x"71"),
  1280 => (x"cb",x"4b",x"74",x"1e"),
  1281 => (x"d8",x"e8",x"c1",x"93"),
  1282 => (x"4a",x"a3",x"c4",x"83"),
  1283 => (x"f2",x"fe",x"49",x"6a"),
  1284 => (x"ca",x"c1",x"87",x"e6"),
  1285 => (x"a3",x"c8",x"7b",x"c3"),
  1286 => (x"51",x"66",x"d4",x"49"),
  1287 => (x"d8",x"49",x"a3",x"c9"),
  1288 => (x"a3",x"ca",x"51",x"66"),
  1289 => (x"51",x"66",x"dc",x"49"),
  1290 => (x"87",x"f5",x"ee",x"26"),
  1291 => (x"5c",x"5b",x"5e",x"0e"),
  1292 => (x"d0",x"ff",x"0e",x"5d"),
  1293 => (x"59",x"a6",x"d8",x"86"),
  1294 => (x"c0",x"48",x"a6",x"c8"),
  1295 => (x"c1",x"80",x"fc",x"78"),
  1296 => (x"c8",x"78",x"66",x"c4"),
  1297 => (x"c4",x"78",x"c1",x"80"),
  1298 => (x"c3",x"78",x"c1",x"80"),
  1299 => (x"c1",x"48",x"ec",x"c2"),
  1300 => (x"d0",x"c2",x"c3",x"78"),
  1301 => (x"48",x"6e",x"7e",x"bf"),
  1302 => (x"cb",x"05",x"a8",x"de"),
  1303 => (x"87",x"d5",x"f3",x"87"),
  1304 => (x"a6",x"cc",x"49",x"70"),
  1305 => (x"87",x"ec",x"d0",x"59"),
  1306 => (x"a8",x"df",x"48",x"6e"),
  1307 => (x"87",x"ee",x"c1",x"05"),
  1308 => (x"49",x"66",x"c0",x"c1"),
  1309 => (x"7e",x"69",x"81",x"c4"),
  1310 => (x"48",x"c9",x"e3",x"c1"),
  1311 => (x"a1",x"d0",x"49",x"6e"),
  1312 => (x"71",x"41",x"20",x"4a"),
  1313 => (x"87",x"f9",x"05",x"aa"),
  1314 => (x"4a",x"c3",x"ca",x"c1"),
  1315 => (x"0a",x"66",x"c0",x"c1"),
  1316 => (x"c0",x"c1",x"0a",x"7a"),
  1317 => (x"81",x"c9",x"49",x"66"),
  1318 => (x"c0",x"c1",x"51",x"df"),
  1319 => (x"81",x"ca",x"49",x"66"),
  1320 => (x"c1",x"51",x"d3",x"c1"),
  1321 => (x"cb",x"49",x"66",x"c0"),
  1322 => (x"4b",x"a1",x"c4",x"81"),
  1323 => (x"6b",x"48",x"a6",x"c4"),
  1324 => (x"72",x"1e",x"71",x"78"),
  1325 => (x"d9",x"e3",x"c1",x"1e"),
  1326 => (x"49",x"66",x"cc",x"48"),
  1327 => (x"20",x"4a",x"a1",x"d0"),
  1328 => (x"05",x"aa",x"71",x"41"),
  1329 => (x"4a",x"26",x"87",x"f9"),
  1330 => (x"79",x"72",x"49",x"26"),
  1331 => (x"df",x"4a",x"a1",x"c9"),
  1332 => (x"c1",x"81",x"ca",x"52"),
  1333 => (x"a6",x"c8",x"51",x"d4"),
  1334 => (x"ce",x"78",x"c2",x"48"),
  1335 => (x"c0",x"e0",x"87",x"f6"),
  1336 => (x"87",x"e2",x"e0",x"87"),
  1337 => (x"87",x"ee",x"df",x"ff"),
  1338 => (x"fb",x"c0",x"4c",x"70"),
  1339 => (x"d2",x"c1",x"02",x"ac"),
  1340 => (x"05",x"66",x"d4",x"87"),
  1341 => (x"c0",x"87",x"c3",x"c1"),
  1342 => (x"1e",x"c1",x"1e",x"1e"),
  1343 => (x"1e",x"cb",x"ea",x"c1"),
  1344 => (x"f2",x"fb",x"49",x"c0"),
  1345 => (x"66",x"d0",x"c1",x"87"),
  1346 => (x"6a",x"82",x"c4",x"4a"),
  1347 => (x"74",x"81",x"c7",x"49"),
  1348 => (x"d8",x"1e",x"c1",x"51"),
  1349 => (x"c8",x"49",x"6a",x"1e"),
  1350 => (x"fd",x"df",x"ff",x"81"),
  1351 => (x"c1",x"86",x"d8",x"87"),
  1352 => (x"c0",x"48",x"66",x"c4"),
  1353 => (x"87",x"c7",x"01",x"a8"),
  1354 => (x"c1",x"48",x"a6",x"c8"),
  1355 => (x"c1",x"87",x"cf",x"78"),
  1356 => (x"c1",x"48",x"66",x"c4"),
  1357 => (x"58",x"a6",x"c8",x"88"),
  1358 => (x"df",x"ff",x"87",x"c4"),
  1359 => (x"a6",x"cc",x"87",x"c8"),
  1360 => (x"74",x"78",x"c2",x"48"),
  1361 => (x"c7",x"cd",x"02",x"9c"),
  1362 => (x"48",x"66",x"c8",x"87"),
  1363 => (x"a8",x"66",x"c8",x"c1"),
  1364 => (x"87",x"fc",x"cc",x"03"),
  1365 => (x"c0",x"48",x"a6",x"d8"),
  1366 => (x"c0",x"80",x"c4",x"78"),
  1367 => (x"f5",x"dd",x"ff",x"78"),
  1368 => (x"c1",x"4c",x"70",x"87"),
  1369 => (x"c2",x"05",x"ac",x"d0"),
  1370 => (x"66",x"dc",x"87",x"db"),
  1371 => (x"87",x"d9",x"e0",x"7e"),
  1372 => (x"e0",x"c0",x"49",x"70"),
  1373 => (x"dd",x"ff",x"59",x"a6"),
  1374 => (x"4c",x"70",x"87",x"dc"),
  1375 => (x"05",x"ac",x"ec",x"c0"),
  1376 => (x"c8",x"87",x"ed",x"c1"),
  1377 => (x"91",x"cb",x"49",x"66"),
  1378 => (x"81",x"66",x"c0",x"c1"),
  1379 => (x"6a",x"4a",x"a1",x"c4"),
  1380 => (x"4a",x"a1",x"c8",x"4d"),
  1381 => (x"c1",x"52",x"66",x"dc"),
  1382 => (x"ff",x"79",x"c4",x"cb"),
  1383 => (x"70",x"87",x"f7",x"dc"),
  1384 => (x"d9",x"02",x"9c",x"4c"),
  1385 => (x"ac",x"fb",x"c0",x"87"),
  1386 => (x"74",x"87",x"d3",x"02"),
  1387 => (x"e5",x"dc",x"ff",x"55"),
  1388 => (x"9c",x"4c",x"70",x"87"),
  1389 => (x"c0",x"87",x"c7",x"02"),
  1390 => (x"ff",x"05",x"ac",x"fb"),
  1391 => (x"e0",x"c0",x"87",x"ed"),
  1392 => (x"55",x"c1",x"c2",x"55"),
  1393 => (x"d4",x"7d",x"97",x"c0"),
  1394 => (x"a9",x"6e",x"49",x"66"),
  1395 => (x"c8",x"87",x"db",x"05"),
  1396 => (x"66",x"c4",x"48",x"66"),
  1397 => (x"87",x"ca",x"04",x"a8"),
  1398 => (x"c1",x"48",x"66",x"c8"),
  1399 => (x"58",x"a6",x"cc",x"80"),
  1400 => (x"66",x"c4",x"87",x"c8"),
  1401 => (x"c8",x"88",x"c1",x"48"),
  1402 => (x"db",x"ff",x"58",x"a6"),
  1403 => (x"4c",x"70",x"87",x"e8"),
  1404 => (x"05",x"ac",x"d0",x"c1"),
  1405 => (x"66",x"d0",x"87",x"c8"),
  1406 => (x"d4",x"80",x"c1",x"48"),
  1407 => (x"d0",x"c1",x"58",x"a6"),
  1408 => (x"e5",x"fd",x"02",x"ac"),
  1409 => (x"a6",x"e0",x"c0",x"87"),
  1410 => (x"78",x"66",x"d4",x"48"),
  1411 => (x"c0",x"48",x"66",x"dc"),
  1412 => (x"05",x"a8",x"66",x"e0"),
  1413 => (x"c0",x"87",x"cb",x"c9"),
  1414 => (x"c0",x"48",x"a6",x"e4"),
  1415 => (x"48",x"74",x"7e",x"78"),
  1416 => (x"c0",x"88",x"fb",x"c0"),
  1417 => (x"70",x"58",x"a6",x"ec"),
  1418 => (x"d0",x"c8",x"02",x"98"),
  1419 => (x"88",x"cb",x"48",x"87"),
  1420 => (x"58",x"a6",x"ec",x"c0"),
  1421 => (x"c1",x"02",x"98",x"70"),
  1422 => (x"c9",x"48",x"87",x"d3"),
  1423 => (x"a6",x"ec",x"c0",x"88"),
  1424 => (x"02",x"98",x"70",x"58"),
  1425 => (x"48",x"87",x"dd",x"c3"),
  1426 => (x"ec",x"c0",x"88",x"c4"),
  1427 => (x"98",x"70",x"58",x"a6"),
  1428 => (x"48",x"87",x"d0",x"02"),
  1429 => (x"ec",x"c0",x"88",x"c1"),
  1430 => (x"98",x"70",x"58",x"a6"),
  1431 => (x"87",x"c4",x"c3",x"02"),
  1432 => (x"d8",x"87",x"d4",x"c7"),
  1433 => (x"f0",x"c0",x"48",x"a6"),
  1434 => (x"e9",x"d9",x"ff",x"78"),
  1435 => (x"c0",x"4c",x"70",x"87"),
  1436 => (x"c0",x"02",x"ac",x"ec"),
  1437 => (x"a6",x"dc",x"87",x"c3"),
  1438 => (x"ac",x"ec",x"c0",x"5c"),
  1439 => (x"87",x"cd",x"c0",x"02"),
  1440 => (x"87",x"d2",x"d9",x"ff"),
  1441 => (x"ec",x"c0",x"4c",x"70"),
  1442 => (x"f3",x"ff",x"05",x"ac"),
  1443 => (x"ac",x"ec",x"c0",x"87"),
  1444 => (x"87",x"c4",x"c0",x"02"),
  1445 => (x"87",x"fe",x"d8",x"ff"),
  1446 => (x"d4",x"1e",x"66",x"d8"),
  1447 => (x"d4",x"1e",x"49",x"66"),
  1448 => (x"c1",x"1e",x"49",x"66"),
  1449 => (x"d8",x"1e",x"cb",x"ea"),
  1450 => (x"ca",x"f5",x"49",x"66"),
  1451 => (x"ca",x"1e",x"c0",x"87"),
  1452 => (x"66",x"e0",x"c0",x"1e"),
  1453 => (x"c1",x"91",x"cb",x"49"),
  1454 => (x"d8",x"81",x"66",x"d8"),
  1455 => (x"a1",x"c4",x"48",x"a6"),
  1456 => (x"bf",x"66",x"d8",x"78"),
  1457 => (x"d1",x"d9",x"ff",x"49"),
  1458 => (x"c0",x"86",x"d8",x"87"),
  1459 => (x"c1",x"06",x"a8",x"b7"),
  1460 => (x"1e",x"c1",x"87",x"c5"),
  1461 => (x"66",x"c8",x"1e",x"de"),
  1462 => (x"d8",x"ff",x"49",x"bf"),
  1463 => (x"86",x"c8",x"87",x"fc"),
  1464 => (x"c0",x"48",x"49",x"70"),
  1465 => (x"a6",x"dc",x"88",x"08"),
  1466 => (x"a8",x"b7",x"c0",x"58"),
  1467 => (x"87",x"e7",x"c0",x"06"),
  1468 => (x"dd",x"48",x"66",x"d8"),
  1469 => (x"de",x"03",x"a8",x"b7"),
  1470 => (x"49",x"bf",x"6e",x"87"),
  1471 => (x"c0",x"81",x"66",x"d8"),
  1472 => (x"66",x"d8",x"51",x"e0"),
  1473 => (x"6e",x"81",x"c1",x"49"),
  1474 => (x"c1",x"c2",x"81",x"bf"),
  1475 => (x"49",x"66",x"d8",x"51"),
  1476 => (x"bf",x"6e",x"81",x"c2"),
  1477 => (x"cc",x"51",x"c0",x"81"),
  1478 => (x"80",x"c1",x"48",x"66"),
  1479 => (x"c1",x"58",x"a6",x"d0"),
  1480 => (x"87",x"d9",x"c4",x"7e"),
  1481 => (x"87",x"e1",x"d9",x"ff"),
  1482 => (x"ff",x"58",x"a6",x"dc"),
  1483 => (x"c0",x"87",x"da",x"d9"),
  1484 => (x"c0",x"58",x"a6",x"ec"),
  1485 => (x"c0",x"05",x"a8",x"ec"),
  1486 => (x"e8",x"c0",x"87",x"ca"),
  1487 => (x"66",x"d8",x"48",x"a6"),
  1488 => (x"87",x"c4",x"c0",x"78"),
  1489 => (x"87",x"ce",x"d6",x"ff"),
  1490 => (x"cb",x"49",x"66",x"c8"),
  1491 => (x"66",x"c0",x"c1",x"91"),
  1492 => (x"70",x"80",x"71",x"48"),
  1493 => (x"c8",x"49",x"6e",x"7e"),
  1494 => (x"ca",x"4a",x"6e",x"81"),
  1495 => (x"52",x"66",x"d8",x"82"),
  1496 => (x"4a",x"66",x"e8",x"c0"),
  1497 => (x"66",x"d8",x"82",x"c1"),
  1498 => (x"72",x"48",x"c1",x"8a"),
  1499 => (x"c1",x"4a",x"70",x"30"),
  1500 => (x"79",x"97",x"72",x"8a"),
  1501 => (x"1e",x"49",x"69",x"97"),
  1502 => (x"c0",x"49",x"66",x"dc"),
  1503 => (x"c4",x"87",x"fc",x"e6"),
  1504 => (x"a6",x"f0",x"c0",x"86"),
  1505 => (x"c4",x"49",x"6e",x"58"),
  1506 => (x"c0",x"4d",x"69",x"81"),
  1507 => (x"dc",x"48",x"66",x"e0"),
  1508 => (x"c0",x"02",x"a8",x"66"),
  1509 => (x"a6",x"d8",x"87",x"c8"),
  1510 => (x"c0",x"78",x"c0",x"48"),
  1511 => (x"a6",x"d8",x"87",x"c5"),
  1512 => (x"d8",x"78",x"c1",x"48"),
  1513 => (x"e0",x"c0",x"1e",x"66"),
  1514 => (x"ff",x"49",x"75",x"1e"),
  1515 => (x"c8",x"87",x"eb",x"d5"),
  1516 => (x"c0",x"4c",x"70",x"86"),
  1517 => (x"c1",x"06",x"ac",x"b7"),
  1518 => (x"85",x"74",x"87",x"d4"),
  1519 => (x"74",x"49",x"e0",x"c0"),
  1520 => (x"c1",x"4b",x"75",x"89"),
  1521 => (x"71",x"4a",x"e9",x"e3"),
  1522 => (x"87",x"dc",x"e3",x"fe"),
  1523 => (x"e4",x"c0",x"85",x"c2"),
  1524 => (x"80",x"c1",x"48",x"66"),
  1525 => (x"58",x"a6",x"e8",x"c0"),
  1526 => (x"49",x"66",x"ec",x"c0"),
  1527 => (x"a9",x"70",x"81",x"c1"),
  1528 => (x"87",x"c8",x"c0",x"02"),
  1529 => (x"c0",x"48",x"a6",x"d8"),
  1530 => (x"87",x"c5",x"c0",x"78"),
  1531 => (x"c1",x"48",x"a6",x"d8"),
  1532 => (x"1e",x"66",x"d8",x"78"),
  1533 => (x"c0",x"49",x"a4",x"c2"),
  1534 => (x"88",x"71",x"48",x"e0"),
  1535 => (x"75",x"1e",x"49",x"70"),
  1536 => (x"d5",x"d4",x"ff",x"49"),
  1537 => (x"c0",x"86",x"c8",x"87"),
  1538 => (x"ff",x"01",x"a8",x"b7"),
  1539 => (x"e4",x"c0",x"87",x"c0"),
  1540 => (x"d1",x"c0",x"02",x"66"),
  1541 => (x"c9",x"49",x"6e",x"87"),
  1542 => (x"66",x"e4",x"c0",x"81"),
  1543 => (x"c1",x"48",x"6e",x"51"),
  1544 => (x"c0",x"78",x"d4",x"cc"),
  1545 => (x"49",x"6e",x"87",x"cc"),
  1546 => (x"51",x"c2",x"81",x"c9"),
  1547 => (x"cd",x"c1",x"48",x"6e"),
  1548 => (x"7e",x"c1",x"78",x"c8"),
  1549 => (x"ff",x"87",x"c6",x"c0"),
  1550 => (x"70",x"87",x"cb",x"d3"),
  1551 => (x"c0",x"02",x"6e",x"4c"),
  1552 => (x"66",x"c8",x"87",x"f5"),
  1553 => (x"a8",x"66",x"c4",x"48"),
  1554 => (x"87",x"cb",x"c0",x"04"),
  1555 => (x"c1",x"48",x"66",x"c8"),
  1556 => (x"58",x"a6",x"cc",x"80"),
  1557 => (x"c4",x"87",x"e0",x"c0"),
  1558 => (x"88",x"c1",x"48",x"66"),
  1559 => (x"c0",x"58",x"a6",x"c8"),
  1560 => (x"c6",x"c1",x"87",x"d5"),
  1561 => (x"c8",x"c0",x"05",x"ac"),
  1562 => (x"48",x"66",x"cc",x"87"),
  1563 => (x"a6",x"d0",x"80",x"c1"),
  1564 => (x"d1",x"d2",x"ff",x"58"),
  1565 => (x"d0",x"4c",x"70",x"87"),
  1566 => (x"80",x"c1",x"48",x"66"),
  1567 => (x"74",x"58",x"a6",x"d4"),
  1568 => (x"cb",x"c0",x"02",x"9c"),
  1569 => (x"48",x"66",x"c8",x"87"),
  1570 => (x"a8",x"66",x"c8",x"c1"),
  1571 => (x"87",x"c4",x"f3",x"04"),
  1572 => (x"87",x"e9",x"d1",x"ff"),
  1573 => (x"c7",x"48",x"66",x"c8"),
  1574 => (x"e5",x"c0",x"03",x"a8"),
  1575 => (x"ec",x"c2",x"c3",x"87"),
  1576 => (x"c8",x"78",x"c0",x"48"),
  1577 => (x"91",x"cb",x"49",x"66"),
  1578 => (x"81",x"66",x"c0",x"c1"),
  1579 => (x"6a",x"4a",x"a1",x"c4"),
  1580 => (x"79",x"52",x"c0",x"4a"),
  1581 => (x"c1",x"48",x"66",x"c8"),
  1582 => (x"58",x"a6",x"cc",x"80"),
  1583 => (x"ff",x"04",x"a8",x"c7"),
  1584 => (x"d0",x"ff",x"87",x"db"),
  1585 => (x"d6",x"dc",x"ff",x"8e"),
  1586 => (x"61",x"6f",x"4c",x"87"),
  1587 => (x"65",x"53",x"20",x"64"),
  1588 => (x"6e",x"69",x"74",x"74"),
  1589 => (x"81",x"20",x"73",x"67"),
  1590 => (x"76",x"61",x"53",x"00"),
  1591 => (x"65",x"53",x"20",x"65"),
  1592 => (x"6e",x"69",x"74",x"74"),
  1593 => (x"81",x"20",x"73",x"67"),
  1594 => (x"00",x"20",x"3a",x"00"),
  1595 => (x"71",x"1e",x"73",x"1e"),
  1596 => (x"c6",x"02",x"9b",x"4b"),
  1597 => (x"e8",x"c2",x"c3",x"87"),
  1598 => (x"c7",x"78",x"c0",x"48"),
  1599 => (x"e8",x"c2",x"c3",x"1e"),
  1600 => (x"c1",x"1e",x"49",x"bf"),
  1601 => (x"c3",x"1e",x"d8",x"e8"),
  1602 => (x"49",x"bf",x"d0",x"c2"),
  1603 => (x"cc",x"87",x"dd",x"ec"),
  1604 => (x"d0",x"c2",x"c3",x"86"),
  1605 => (x"d3",x"e7",x"49",x"bf"),
  1606 => (x"02",x"9b",x"73",x"87"),
  1607 => (x"e8",x"c1",x"87",x"c8"),
  1608 => (x"f6",x"c0",x"49",x"d8"),
  1609 => (x"da",x"ff",x"87",x"f9"),
  1610 => (x"c1",x"1e",x"87",x"f9"),
  1611 => (x"c1",x"49",x"c6",x"e5"),
  1612 => (x"c1",x"87",x"cf",x"ce"),
  1613 => (x"c0",x"48",x"e5",x"e7"),
  1614 => (x"fb",x"e9",x"c1",x"50"),
  1615 => (x"d6",x"ff",x"49",x"bf"),
  1616 => (x"48",x"c0",x"87",x"e5"),
  1617 => (x"4f",x"43",x"4f",x"26"),
  1618 => (x"20",x"20",x"45",x"52"),
  1619 => (x"46",x"43",x"20",x"20"),
  1620 => (x"ce",x"1e",x"00",x"47"),
  1621 => (x"49",x"c1",x"87",x"c8"),
  1622 => (x"fe",x"87",x"d1",x"fe"),
  1623 => (x"70",x"87",x"fe",x"e5"),
  1624 => (x"87",x"cd",x"02",x"98"),
  1625 => (x"87",x"f9",x"ee",x"fe"),
  1626 => (x"c4",x"02",x"98",x"70"),
  1627 => (x"c2",x"4a",x"c1",x"87"),
  1628 => (x"72",x"4a",x"c0",x"87"),
  1629 => (x"87",x"ce",x"05",x"9a"),
  1630 => (x"e6",x"c1",x"1e",x"c0"),
  1631 => (x"c1",x"c1",x"49",x"e6"),
  1632 => (x"86",x"c4",x"87",x"fa"),
  1633 => (x"cb",x"c1",x"87",x"fe"),
  1634 => (x"1e",x"c0",x"87",x"e2"),
  1635 => (x"49",x"f1",x"e6",x"c1"),
  1636 => (x"87",x"e8",x"c1",x"c1"),
  1637 => (x"d1",x"fe",x"1e",x"c0"),
  1638 => (x"c1",x"49",x"70",x"87"),
  1639 => (x"c4",x"87",x"dd",x"c1"),
  1640 => (x"8e",x"f8",x"87",x"c7"),
  1641 => (x"44",x"53",x"4f",x"26"),
  1642 => (x"69",x"61",x"66",x"20"),
  1643 => (x"2e",x"64",x"65",x"6c"),
  1644 => (x"6f",x"6f",x"42",x"00"),
  1645 => (x"67",x"6e",x"69",x"74"),
  1646 => (x"00",x"2e",x"2e",x"2e"),
  1647 => (x"d4",x"49",x"c0",x"1e"),
  1648 => (x"f8",x"c0",x"87",x"e2"),
  1649 => (x"c4",x"c1",x"87",x"f9"),
  1650 => (x"87",x"f1",x"87",x"e8"),
  1651 => (x"c3",x"1e",x"4f",x"26"),
  1652 => (x"c0",x"48",x"e8",x"c2"),
  1653 => (x"d0",x"c2",x"c3",x"78"),
  1654 => (x"fd",x"78",x"c0",x"48"),
  1655 => (x"db",x"ff",x"87",x"f4"),
  1656 => (x"26",x"48",x"c0",x"87"),
  1657 => (x"20",x"00",x"00",x"4f"),
  1658 => (x"20",x"20",x"20",x"20"),
  1659 => (x"20",x"20",x"20",x"20"),
  1660 => (x"20",x"20",x"20",x"20"),
  1661 => (x"74",x"69",x"78",x"45"),
  1662 => (x"20",x"20",x"20",x"20"),
  1663 => (x"20",x"20",x"20",x"20"),
  1664 => (x"20",x"20",x"20",x"20"),
  1665 => (x"20",x"80",x"00",x"81"),
  1666 => (x"20",x"20",x"20",x"20"),
  1667 => (x"20",x"20",x"20",x"20"),
  1668 => (x"42",x"20",x"20",x"20"),
  1669 => (x"00",x"6b",x"63",x"61"),
  1670 => (x"00",x"00",x"12",x"c4"),
  1671 => (x"00",x"00",x"30",x"bc"),
  1672 => (x"c4",x"00",x"00",x"00"),
  1673 => (x"da",x"00",x"00",x"12"),
  1674 => (x"00",x"00",x"00",x"30"),
  1675 => (x"12",x"c4",x"00",x"00"),
  1676 => (x"30",x"f8",x"00",x"00"),
  1677 => (x"00",x"00",x"00",x"00"),
  1678 => (x"00",x"12",x"c4",x"00"),
  1679 => (x"00",x"31",x"16",x"00"),
  1680 => (x"00",x"00",x"00",x"00"),
  1681 => (x"00",x"00",x"12",x"c4"),
  1682 => (x"00",x"00",x"31",x"34"),
  1683 => (x"c4",x"00",x"00",x"00"),
  1684 => (x"52",x"00",x"00",x"12"),
  1685 => (x"00",x"00",x"00",x"31"),
  1686 => (x"12",x"c4",x"00",x"00"),
  1687 => (x"31",x"70",x"00",x"00"),
  1688 => (x"00",x"00",x"00",x"00"),
  1689 => (x"00",x"12",x"c4",x"00"),
  1690 => (x"00",x"00",x"00",x"00"),
  1691 => (x"00",x"00",x"00",x"00"),
  1692 => (x"00",x"00",x"13",x"59"),
  1693 => (x"00",x"00",x"00",x"00"),
  1694 => (x"7f",x"00",x"00",x"00"),
  1695 => (x"43",x"00",x"00",x"1a"),
  1696 => (x"20",x"20",x"34",x"36"),
  1697 => (x"52",x"20",x"20",x"20"),
  1698 => (x"4c",x"00",x"4d",x"4f"),
  1699 => (x"20",x"64",x"61",x"6f"),
  1700 => (x"1e",x"00",x"2e",x"2a"),
  1701 => (x"c0",x"48",x"f0",x"fe"),
  1702 => (x"79",x"09",x"cd",x"78"),
  1703 => (x"1e",x"4f",x"26",x"09"),
  1704 => (x"bf",x"f0",x"fe",x"1e"),
  1705 => (x"26",x"26",x"48",x"7e"),
  1706 => (x"f0",x"fe",x"1e",x"4f"),
  1707 => (x"26",x"78",x"c1",x"48"),
  1708 => (x"f0",x"fe",x"1e",x"4f"),
  1709 => (x"26",x"78",x"c0",x"48"),
  1710 => (x"4a",x"71",x"1e",x"4f"),
  1711 => (x"c1",x"7a",x"97",x"c0"),
  1712 => (x"51",x"c0",x"49",x"a2"),
  1713 => (x"c0",x"49",x"a2",x"ca"),
  1714 => (x"49",x"a2",x"cb",x"51"),
  1715 => (x"4f",x"26",x"51",x"c0"),
  1716 => (x"5c",x"5b",x"5e",x"0e"),
  1717 => (x"71",x"86",x"f0",x"0e"),
  1718 => (x"49",x"a4",x"ca",x"4c"),
  1719 => (x"cb",x"7e",x"69",x"97"),
  1720 => (x"6b",x"97",x"4b",x"a4"),
  1721 => (x"58",x"a6",x"c8",x"48"),
  1722 => (x"a6",x"cc",x"80",x"c1"),
  1723 => (x"d0",x"98",x"c7",x"58"),
  1724 => (x"48",x"6e",x"58",x"a6"),
  1725 => (x"05",x"a8",x"66",x"cc"),
  1726 => (x"69",x"97",x"87",x"db"),
  1727 => (x"48",x"6b",x"97",x"7e"),
  1728 => (x"c1",x"58",x"a6",x"c8"),
  1729 => (x"58",x"a6",x"cc",x"80"),
  1730 => (x"a6",x"d0",x"98",x"c7"),
  1731 => (x"cc",x"48",x"6e",x"58"),
  1732 => (x"e5",x"02",x"a8",x"66"),
  1733 => (x"87",x"d9",x"fe",x"87"),
  1734 => (x"97",x"4a",x"a4",x"cc"),
  1735 => (x"a1",x"72",x"49",x"6b"),
  1736 => (x"51",x"66",x"dc",x"49"),
  1737 => (x"6e",x"7e",x"6b",x"97"),
  1738 => (x"c8",x"80",x"c1",x"48"),
  1739 => (x"98",x"c7",x"58",x"a6"),
  1740 => (x"70",x"58",x"a6",x"cc"),
  1741 => (x"d2",x"c3",x"7b",x"97"),
  1742 => (x"87",x"ed",x"fd",x"87"),
  1743 => (x"87",x"c2",x"8e",x"f0"),
  1744 => (x"4c",x"26",x"4d",x"26"),
  1745 => (x"4f",x"26",x"4b",x"26"),
  1746 => (x"5c",x"5b",x"5e",x"0e"),
  1747 => (x"86",x"f4",x"0e",x"5d"),
  1748 => (x"6d",x"97",x"4d",x"71"),
  1749 => (x"4c",x"a5",x"c1",x"7e"),
  1750 => (x"c8",x"48",x"6c",x"97"),
  1751 => (x"48",x"6e",x"58",x"a6"),
  1752 => (x"05",x"a8",x"66",x"c4"),
  1753 => (x"48",x"ff",x"87",x"c5"),
  1754 => (x"fd",x"87",x"e6",x"c0"),
  1755 => (x"a5",x"c2",x"87",x"c3"),
  1756 => (x"4b",x"6c",x"97",x"49"),
  1757 => (x"97",x"4b",x"a3",x"71"),
  1758 => (x"6c",x"97",x"4b",x"6b"),
  1759 => (x"c1",x"48",x"6e",x"7e"),
  1760 => (x"58",x"a6",x"c8",x"80"),
  1761 => (x"a6",x"cc",x"98",x"c7"),
  1762 => (x"7c",x"97",x"70",x"58"),
  1763 => (x"73",x"87",x"da",x"fc"),
  1764 => (x"fe",x"8e",x"f4",x"48"),
  1765 => (x"5e",x"0e",x"87",x"ea"),
  1766 => (x"f4",x"0e",x"5c",x"5b"),
  1767 => (x"d8",x"4c",x"71",x"86"),
  1768 => (x"ff",x"c3",x"4a",x"66"),
  1769 => (x"4b",x"a4",x"c2",x"9a"),
  1770 => (x"73",x"49",x"6c",x"97"),
  1771 => (x"51",x"72",x"49",x"a1"),
  1772 => (x"6e",x"7e",x"6c",x"97"),
  1773 => (x"c8",x"80",x"c1",x"48"),
  1774 => (x"98",x"c7",x"58",x"a6"),
  1775 => (x"70",x"58",x"a6",x"cc"),
  1776 => (x"fd",x"8e",x"f4",x"54"),
  1777 => (x"f0",x"1e",x"87",x"fc"),
  1778 => (x"7e",x"69",x"97",x"86"),
  1779 => (x"97",x"4a",x"a1",x"c1"),
  1780 => (x"a6",x"c8",x"48",x"6a"),
  1781 => (x"c4",x"48",x"6e",x"58"),
  1782 => (x"04",x"a8",x"b7",x"66"),
  1783 => (x"69",x"97",x"87",x"d3"),
  1784 => (x"48",x"6a",x"97",x"7e"),
  1785 => (x"6e",x"58",x"a6",x"c8"),
  1786 => (x"88",x"66",x"c4",x"48"),
  1787 => (x"d6",x"58",x"a6",x"cc"),
  1788 => (x"6e",x"7e",x"11",x"87"),
  1789 => (x"a6",x"80",x"c8",x"48"),
  1790 => (x"cc",x"48",x"12",x"58"),
  1791 => (x"66",x"c4",x"58",x"a6"),
  1792 => (x"88",x"66",x"c8",x"48"),
  1793 => (x"f0",x"58",x"a6",x"d0"),
  1794 => (x"1e",x"4f",x"26",x"8e"),
  1795 => (x"86",x"f4",x"1e",x"73"),
  1796 => (x"e0",x"87",x"de",x"fa"),
  1797 => (x"c0",x"49",x"4b",x"bf"),
  1798 => (x"02",x"99",x"c0",x"e0"),
  1799 => (x"1e",x"73",x"87",x"cb"),
  1800 => (x"49",x"ce",x"c6",x"c3"),
  1801 => (x"c4",x"87",x"ef",x"fd"),
  1802 => (x"d0",x"49",x"73",x"86"),
  1803 => (x"c1",x"02",x"99",x"c0"),
  1804 => (x"c6",x"c3",x"87",x"c0"),
  1805 => (x"7e",x"bf",x"97",x"d8"),
  1806 => (x"97",x"d9",x"c6",x"c3"),
  1807 => (x"a6",x"c8",x"48",x"bf"),
  1808 => (x"c4",x"48",x"6e",x"58"),
  1809 => (x"c0",x"02",x"a8",x"66"),
  1810 => (x"c6",x"c3",x"87",x"e8"),
  1811 => (x"49",x"bf",x"97",x"d8"),
  1812 => (x"81",x"da",x"c6",x"c3"),
  1813 => (x"08",x"e0",x"48",x"11"),
  1814 => (x"d8",x"c6",x"c3",x"78"),
  1815 => (x"6e",x"7e",x"bf",x"97"),
  1816 => (x"c8",x"80",x"c1",x"48"),
  1817 => (x"98",x"c7",x"58",x"a6"),
  1818 => (x"c3",x"58",x"a6",x"cc"),
  1819 => (x"c8",x"48",x"d8",x"c6"),
  1820 => (x"bf",x"e4",x"50",x"66"),
  1821 => (x"e0",x"c0",x"49",x"4b"),
  1822 => (x"cb",x"02",x"99",x"c0"),
  1823 => (x"c3",x"1e",x"73",x"87"),
  1824 => (x"fc",x"49",x"e2",x"c6"),
  1825 => (x"86",x"c4",x"87",x"d0"),
  1826 => (x"c0",x"d0",x"49",x"73"),
  1827 => (x"c0",x"c1",x"02",x"99"),
  1828 => (x"ec",x"c6",x"c3",x"87"),
  1829 => (x"c3",x"7e",x"bf",x"97"),
  1830 => (x"bf",x"97",x"ed",x"c6"),
  1831 => (x"58",x"a6",x"c8",x"48"),
  1832 => (x"66",x"c4",x"48",x"6e"),
  1833 => (x"e8",x"c0",x"02",x"a8"),
  1834 => (x"ec",x"c6",x"c3",x"87"),
  1835 => (x"c3",x"49",x"bf",x"97"),
  1836 => (x"11",x"81",x"ee",x"c6"),
  1837 => (x"78",x"08",x"e4",x"48"),
  1838 => (x"97",x"ec",x"c6",x"c3"),
  1839 => (x"48",x"6e",x"7e",x"bf"),
  1840 => (x"a6",x"c8",x"80",x"c1"),
  1841 => (x"cc",x"98",x"c7",x"58"),
  1842 => (x"c6",x"c3",x"58",x"a6"),
  1843 => (x"66",x"c8",x"48",x"ec"),
  1844 => (x"87",x"cb",x"f7",x"50"),
  1845 => (x"d0",x"f7",x"7e",x"70"),
  1846 => (x"f9",x"8e",x"f4",x"87"),
  1847 => (x"c3",x"1e",x"87",x"e6"),
  1848 => (x"f7",x"49",x"ce",x"c6"),
  1849 => (x"c6",x"c3",x"87",x"d3"),
  1850 => (x"cc",x"f7",x"49",x"e2"),
  1851 => (x"cb",x"f0",x"c1",x"87"),
  1852 => (x"87",x"df",x"f6",x"49"),
  1853 => (x"26",x"87",x"c8",x"c4"),
  1854 => (x"d0",x"ff",x"1e",x"4f"),
  1855 => (x"78",x"e1",x"c8",x"48"),
  1856 => (x"c5",x"48",x"d4",x"ff"),
  1857 => (x"02",x"66",x"c4",x"78"),
  1858 => (x"e0",x"c3",x"87",x"c3"),
  1859 => (x"02",x"66",x"c8",x"78"),
  1860 => (x"d4",x"ff",x"87",x"c6"),
  1861 => (x"78",x"f0",x"c3",x"48"),
  1862 => (x"71",x"48",x"d4",x"ff"),
  1863 => (x"48",x"d0",x"ff",x"78"),
  1864 => (x"c0",x"78",x"e1",x"c8"),
  1865 => (x"4f",x"26",x"78",x"e0"),
  1866 => (x"5c",x"5b",x"5e",x"0e"),
  1867 => (x"c3",x"4c",x"71",x"0e"),
  1868 => (x"f8",x"49",x"ce",x"c6"),
  1869 => (x"4a",x"70",x"87",x"d2"),
  1870 => (x"04",x"aa",x"b7",x"c0"),
  1871 => (x"c3",x"87",x"e3",x"c2"),
  1872 => (x"c9",x"05",x"aa",x"e0"),
  1873 => (x"f2",x"f7",x"c1",x"87"),
  1874 => (x"c2",x"78",x"c1",x"48"),
  1875 => (x"f0",x"c3",x"87",x"d4"),
  1876 => (x"87",x"c9",x"05",x"aa"),
  1877 => (x"48",x"ee",x"f7",x"c1"),
  1878 => (x"f5",x"c1",x"78",x"c1"),
  1879 => (x"f2",x"f7",x"c1",x"87"),
  1880 => (x"87",x"c7",x"02",x"bf"),
  1881 => (x"c0",x"c2",x"4b",x"72"),
  1882 => (x"72",x"87",x"c2",x"b3"),
  1883 => (x"05",x"9c",x"74",x"4b"),
  1884 => (x"f7",x"c1",x"87",x"d1"),
  1885 => (x"c1",x"1e",x"bf",x"ee"),
  1886 => (x"1e",x"bf",x"f2",x"f7"),
  1887 => (x"f8",x"fd",x"49",x"72"),
  1888 => (x"c1",x"86",x"c8",x"87"),
  1889 => (x"02",x"bf",x"ee",x"f7"),
  1890 => (x"73",x"87",x"e0",x"c0"),
  1891 => (x"29",x"b7",x"c4",x"49"),
  1892 => (x"ce",x"f9",x"c1",x"91"),
  1893 => (x"cf",x"4a",x"73",x"81"),
  1894 => (x"c1",x"92",x"c2",x"9a"),
  1895 => (x"70",x"30",x"72",x"48"),
  1896 => (x"72",x"ba",x"ff",x"4a"),
  1897 => (x"70",x"98",x"69",x"48"),
  1898 => (x"73",x"87",x"db",x"79"),
  1899 => (x"29",x"b7",x"c4",x"49"),
  1900 => (x"ce",x"f9",x"c1",x"91"),
  1901 => (x"cf",x"4a",x"73",x"81"),
  1902 => (x"c3",x"92",x"c2",x"9a"),
  1903 => (x"70",x"30",x"72",x"48"),
  1904 => (x"b0",x"69",x"48",x"4a"),
  1905 => (x"f7",x"c1",x"79",x"70"),
  1906 => (x"78",x"c0",x"48",x"f2"),
  1907 => (x"48",x"ee",x"f7",x"c1"),
  1908 => (x"c6",x"c3",x"78",x"c0"),
  1909 => (x"ef",x"f5",x"49",x"ce"),
  1910 => (x"c0",x"4a",x"70",x"87"),
  1911 => (x"fd",x"03",x"aa",x"b7"),
  1912 => (x"48",x"c0",x"87",x"dd"),
  1913 => (x"4d",x"26",x"87",x"c2"),
  1914 => (x"4b",x"26",x"4c",x"26"),
  1915 => (x"00",x"00",x"4f",x"26"),
  1916 => (x"00",x"00",x"00",x"00"),
  1917 => (x"71",x"1e",x"00",x"00"),
  1918 => (x"eb",x"fc",x"49",x"4a"),
  1919 => (x"1e",x"4f",x"26",x"87"),
  1920 => (x"49",x"72",x"4a",x"c0"),
  1921 => (x"f9",x"c1",x"91",x"c4"),
  1922 => (x"79",x"c0",x"81",x"ce"),
  1923 => (x"b7",x"d0",x"82",x"c1"),
  1924 => (x"87",x"ee",x"04",x"aa"),
  1925 => (x"5e",x"0e",x"4f",x"26"),
  1926 => (x"0e",x"5d",x"5c",x"5b"),
  1927 => (x"d0",x"f2",x"4d",x"71"),
  1928 => (x"c4",x"4a",x"75",x"87"),
  1929 => (x"c1",x"92",x"2a",x"b7"),
  1930 => (x"75",x"82",x"ce",x"f9"),
  1931 => (x"c2",x"9c",x"cf",x"4c"),
  1932 => (x"4b",x"49",x"6a",x"94"),
  1933 => (x"9b",x"c3",x"2b",x"74"),
  1934 => (x"30",x"74",x"48",x"c2"),
  1935 => (x"bc",x"ff",x"4c",x"70"),
  1936 => (x"98",x"71",x"48",x"74"),
  1937 => (x"e0",x"f1",x"7a",x"70"),
  1938 => (x"fe",x"48",x"73",x"87"),
  1939 => (x"00",x"00",x"87",x"d8"),
  1940 => (x"00",x"00",x"00",x"00"),
  1941 => (x"00",x"00",x"00",x"00"),
  1942 => (x"00",x"00",x"00",x"00"),
  1943 => (x"00",x"00",x"00",x"00"),
  1944 => (x"00",x"00",x"00",x"00"),
  1945 => (x"00",x"00",x"00",x"00"),
  1946 => (x"00",x"00",x"00",x"00"),
  1947 => (x"00",x"00",x"00",x"00"),
  1948 => (x"00",x"00",x"00",x"00"),
  1949 => (x"00",x"00",x"00",x"00"),
  1950 => (x"00",x"00",x"00",x"00"),
  1951 => (x"00",x"00",x"00",x"00"),
  1952 => (x"00",x"00",x"00",x"00"),
  1953 => (x"00",x"00",x"00",x"00"),
  1954 => (x"00",x"00",x"00",x"00"),
  1955 => (x"73",x"1e",x"00",x"00"),
  1956 => (x"c3",x"4b",x"71",x"1e"),
  1957 => (x"f2",x"49",x"e2",x"c6"),
  1958 => (x"49",x"70",x"87",x"ee"),
  1959 => (x"49",x"f0",x"c1",x"1e"),
  1960 => (x"c4",x"87",x"cb",x"c8"),
  1961 => (x"e2",x"c6",x"c3",x"86"),
  1962 => (x"87",x"dc",x"f2",x"49"),
  1963 => (x"d4",x"ff",x"49",x"70"),
  1964 => (x"c3",x"78",x"71",x"48"),
  1965 => (x"f2",x"49",x"e2",x"c6"),
  1966 => (x"49",x"70",x"87",x"ce"),
  1967 => (x"71",x"48",x"d4",x"ff"),
  1968 => (x"05",x"ab",x"c4",x"78"),
  1969 => (x"c6",x"c3",x"87",x"ce"),
  1970 => (x"fb",x"f1",x"49",x"e2"),
  1971 => (x"ff",x"49",x"70",x"87"),
  1972 => (x"78",x"71",x"48",x"d4"),
  1973 => (x"c0",x"48",x"d0",x"ff"),
  1974 => (x"87",x"c4",x"78",x"e0"),
  1975 => (x"4c",x"26",x"4d",x"26"),
  1976 => (x"4f",x"26",x"4b",x"26"),
  1977 => (x"5c",x"5b",x"5e",x"0e"),
  1978 => (x"4a",x"71",x"0e",x"5d"),
  1979 => (x"87",x"c6",x"02",x"9a"),
  1980 => (x"48",x"ff",x"c1",x"c2"),
  1981 => (x"c1",x"c2",x"78",x"c0"),
  1982 => (x"c1",x"05",x"bf",x"ff"),
  1983 => (x"c6",x"c3",x"87",x"c6"),
  1984 => (x"c3",x"f1",x"49",x"e2"),
  1985 => (x"a8",x"b7",x"c0",x"87"),
  1986 => (x"c3",x"87",x"cd",x"04"),
  1987 => (x"f0",x"49",x"e2",x"c6"),
  1988 => (x"b7",x"c0",x"87",x"f6"),
  1989 => (x"87",x"f3",x"03",x"a8"),
  1990 => (x"bf",x"ff",x"c1",x"c2"),
  1991 => (x"ff",x"c1",x"c2",x"49"),
  1992 => (x"78",x"a1",x"c1",x"48"),
  1993 => (x"81",x"cf",x"c2",x"c2"),
  1994 => (x"c2",x"c2",x"48",x"11"),
  1995 => (x"c2",x"c2",x"58",x"c7"),
  1996 => (x"78",x"c0",x"48",x"c7"),
  1997 => (x"c0",x"49",x"f2",x"c0"),
  1998 => (x"70",x"87",x"de",x"ec"),
  1999 => (x"fa",x"c6",x"c3",x"49"),
  2000 => (x"87",x"f8",x"c4",x"59"),
  2001 => (x"bf",x"c7",x"c2",x"c2"),
  2002 => (x"87",x"f2",x"c1",x"02"),
  2003 => (x"49",x"e2",x"c6",x"c3"),
  2004 => (x"c0",x"87",x"f5",x"ef"),
  2005 => (x"cd",x"04",x"a8",x"b7"),
  2006 => (x"c7",x"c2",x"c2",x"87"),
  2007 => (x"88",x"c1",x"48",x"bf"),
  2008 => (x"58",x"cb",x"c2",x"c2"),
  2009 => (x"c6",x"c3",x"87",x"db"),
  2010 => (x"c0",x"49",x"bf",x"f6"),
  2011 => (x"70",x"87",x"f6",x"eb"),
  2012 => (x"87",x"cd",x"02",x"98"),
  2013 => (x"49",x"e2",x"c6",x"c3"),
  2014 => (x"c2",x"87",x"fe",x"ec"),
  2015 => (x"c0",x"48",x"ff",x"c1"),
  2016 => (x"c3",x"c2",x"c2",x"78"),
  2017 => (x"f3",x"c3",x"05",x"bf"),
  2018 => (x"c7",x"c2",x"c2",x"87"),
  2019 => (x"eb",x"c3",x"05",x"bf"),
  2020 => (x"ff",x"c1",x"c2",x"87"),
  2021 => (x"c1",x"c2",x"49",x"bf"),
  2022 => (x"a1",x"c1",x"48",x"ff"),
  2023 => (x"cf",x"c2",x"c2",x"78"),
  2024 => (x"49",x"4b",x"11",x"81"),
  2025 => (x"02",x"99",x"c0",x"c2"),
  2026 => (x"73",x"87",x"cc",x"c0"),
  2027 => (x"98",x"ff",x"c1",x"48"),
  2028 => (x"58",x"cb",x"c2",x"c2"),
  2029 => (x"c2",x"87",x"c5",x"c3"),
  2030 => (x"c2",x"5b",x"c7",x"c2"),
  2031 => (x"c2",x"c2",x"87",x"fe"),
  2032 => (x"c1",x"02",x"bf",x"c3"),
  2033 => (x"c6",x"c3",x"87",x"db"),
  2034 => (x"c0",x"49",x"bf",x"f6"),
  2035 => (x"70",x"87",x"d6",x"ea"),
  2036 => (x"e7",x"c2",x"02",x"98"),
  2037 => (x"ff",x"c1",x"c2",x"87"),
  2038 => (x"c1",x"c2",x"49",x"bf"),
  2039 => (x"a1",x"c1",x"48",x"ff"),
  2040 => (x"cf",x"c2",x"c2",x"78"),
  2041 => (x"49",x"69",x"97",x"81"),
  2042 => (x"e2",x"c6",x"c3",x"1e"),
  2043 => (x"87",x"e0",x"eb",x"49"),
  2044 => (x"c2",x"c2",x"86",x"c4"),
  2045 => (x"c1",x"49",x"bf",x"c3"),
  2046 => (x"c7",x"c2",x"c2",x"89"),
  2047 => (x"c7",x"c2",x"c2",x"59"),
  2048 => (x"71",x"78",x"c1",x"48"),
  2049 => (x"c6",x"c0",x"02",x"99"),
  2050 => (x"4c",x"f2",x"c0",x"87"),
  2051 => (x"d7",x"87",x"c3",x"c0"),
  2052 => (x"49",x"74",x"4c",x"dc"),
  2053 => (x"87",x"c1",x"e9",x"c0"),
  2054 => (x"c6",x"c3",x"49",x"70"),
  2055 => (x"db",x"c1",x"59",x"fa"),
  2056 => (x"e2",x"c6",x"c3",x"87"),
  2057 => (x"87",x"de",x"ee",x"49"),
  2058 => (x"02",x"9b",x"4b",x"70"),
  2059 => (x"c2",x"87",x"ee",x"c0"),
  2060 => (x"b7",x"bf",x"cb",x"c2"),
  2061 => (x"e4",x"c0",x"03",x"ab"),
  2062 => (x"f6",x"c6",x"c3",x"87"),
  2063 => (x"e8",x"c0",x"49",x"bf"),
  2064 => (x"98",x"70",x"87",x"e3"),
  2065 => (x"87",x"f4",x"c0",x"02"),
  2066 => (x"c2",x"c2",x"48",x"c7"),
  2067 => (x"c2",x"88",x"bf",x"cb"),
  2068 => (x"c3",x"58",x"cf",x"c2"),
  2069 => (x"e9",x"49",x"e2",x"c6"),
  2070 => (x"df",x"c0",x"87",x"df"),
  2071 => (x"49",x"dc",x"d7",x"87"),
  2072 => (x"87",x"f5",x"e7",x"c0"),
  2073 => (x"c6",x"c3",x"49",x"70"),
  2074 => (x"c2",x"c2",x"59",x"fa"),
  2075 => (x"b7",x"4a",x"bf",x"cb"),
  2076 => (x"c7",x"c0",x"04",x"ab"),
  2077 => (x"d5",x"f8",x"49",x"87"),
  2078 => (x"87",x"e5",x"fe",x"87"),
  2079 => (x"00",x"87",x"dd",x"f9"),
  2080 => (x"00",x"00",x"00",x"00"),
  2081 => (x"00",x"00",x"00",x"00"),
  2082 => (x"04",x"00",x"00",x"00"),
  2083 => (x"01",x"00",x"00",x"00"),
  2084 => (x"f3",x"08",x"82",x"ff"),
  2085 => (x"f3",x"64",x"f3",x"c8"),
  2086 => (x"81",x"01",x"f2",x"50"),
  2087 => (x"1e",x"00",x"f4",x"01"),
  2088 => (x"c8",x"48",x"d0",x"ff"),
  2089 => (x"48",x"71",x"78",x"e1"),
  2090 => (x"78",x"08",x"d4",x"ff"),
  2091 => (x"ff",x"1e",x"4f",x"26"),
  2092 => (x"e1",x"c8",x"48",x"d0"),
  2093 => (x"ff",x"48",x"71",x"78"),
  2094 => (x"c4",x"78",x"08",x"d4"),
  2095 => (x"d4",x"ff",x"48",x"66"),
  2096 => (x"4f",x"26",x"78",x"08"),
  2097 => (x"c4",x"4a",x"71",x"1e"),
  2098 => (x"72",x"1e",x"49",x"66"),
  2099 => (x"87",x"de",x"ff",x"49"),
  2100 => (x"c0",x"48",x"d0",x"ff"),
  2101 => (x"26",x"26",x"78",x"e0"),
  2102 => (x"1e",x"73",x"1e",x"4f"),
  2103 => (x"66",x"c8",x"4b",x"71"),
  2104 => (x"4a",x"73",x"1e",x"49"),
  2105 => (x"49",x"a2",x"e0",x"c1"),
  2106 => (x"26",x"87",x"d9",x"ff"),
  2107 => (x"4d",x"26",x"87",x"c4"),
  2108 => (x"4b",x"26",x"4c",x"26"),
  2109 => (x"ff",x"1e",x"4f",x"26"),
  2110 => (x"ff",x"c3",x"4a",x"d4"),
  2111 => (x"48",x"d0",x"ff",x"7a"),
  2112 => (x"de",x"78",x"e1",x"c8"),
  2113 => (x"fa",x"c6",x"c3",x"7a"),
  2114 => (x"48",x"49",x"7a",x"bf"),
  2115 => (x"7a",x"70",x"28",x"c8"),
  2116 => (x"28",x"d0",x"48",x"71"),
  2117 => (x"48",x"71",x"7a",x"70"),
  2118 => (x"7a",x"70",x"28",x"d8"),
  2119 => (x"bf",x"fe",x"c6",x"c3"),
  2120 => (x"c8",x"48",x"49",x"7a"),
  2121 => (x"71",x"7a",x"70",x"28"),
  2122 => (x"70",x"28",x"d0",x"48"),
  2123 => (x"d8",x"48",x"71",x"7a"),
  2124 => (x"ff",x"7a",x"70",x"28"),
  2125 => (x"e0",x"c0",x"48",x"d0"),
  2126 => (x"1e",x"4f",x"26",x"78"),
  2127 => (x"4a",x"71",x"1e",x"73"),
  2128 => (x"bf",x"fa",x"c6",x"c3"),
  2129 => (x"c0",x"2b",x"72",x"4b"),
  2130 => (x"ce",x"04",x"aa",x"e0"),
  2131 => (x"c0",x"49",x"72",x"87"),
  2132 => (x"c6",x"c3",x"89",x"e0"),
  2133 => (x"71",x"4b",x"bf",x"fe"),
  2134 => (x"c0",x"87",x"cf",x"2b"),
  2135 => (x"89",x"72",x"49",x"e0"),
  2136 => (x"bf",x"fe",x"c6",x"c3"),
  2137 => (x"70",x"30",x"71",x"48"),
  2138 => (x"66",x"c8",x"b3",x"49"),
  2139 => (x"c4",x"48",x"73",x"9b"),
  2140 => (x"26",x"4d",x"26",x"87"),
  2141 => (x"26",x"4b",x"26",x"4c"),
  2142 => (x"5b",x"5e",x"0e",x"4f"),
  2143 => (x"ec",x"0e",x"5d",x"5c"),
  2144 => (x"c3",x"4b",x"71",x"86"),
  2145 => (x"7e",x"bf",x"fa",x"c6"),
  2146 => (x"c0",x"2c",x"73",x"4c"),
  2147 => (x"c0",x"04",x"ab",x"e0"),
  2148 => (x"a6",x"c4",x"87",x"e0"),
  2149 => (x"73",x"78",x"c0",x"48"),
  2150 => (x"89",x"e0",x"c0",x"49"),
  2151 => (x"e4",x"c0",x"4a",x"71"),
  2152 => (x"30",x"72",x"48",x"66"),
  2153 => (x"c3",x"58",x"a6",x"cc"),
  2154 => (x"4d",x"bf",x"fe",x"c6"),
  2155 => (x"c0",x"2c",x"71",x"4c"),
  2156 => (x"49",x"73",x"87",x"e4"),
  2157 => (x"48",x"66",x"e4",x"c0"),
  2158 => (x"a6",x"c8",x"30",x"71"),
  2159 => (x"49",x"e0",x"c0",x"58"),
  2160 => (x"e4",x"c0",x"89",x"73"),
  2161 => (x"28",x"71",x"48",x"66"),
  2162 => (x"c3",x"58",x"a6",x"cc"),
  2163 => (x"4d",x"bf",x"fe",x"c6"),
  2164 => (x"70",x"30",x"71",x"48"),
  2165 => (x"e4",x"c0",x"b4",x"49"),
  2166 => (x"84",x"c1",x"9c",x"66"),
  2167 => (x"ac",x"66",x"e8",x"c0"),
  2168 => (x"c0",x"87",x"c2",x"04"),
  2169 => (x"ab",x"e0",x"c0",x"4c"),
  2170 => (x"cc",x"87",x"d3",x"04"),
  2171 => (x"78",x"c0",x"48",x"a6"),
  2172 => (x"e0",x"c0",x"49",x"73"),
  2173 => (x"71",x"48",x"74",x"89"),
  2174 => (x"58",x"a6",x"d4",x"30"),
  2175 => (x"49",x"73",x"87",x"d5"),
  2176 => (x"30",x"71",x"48",x"74"),
  2177 => (x"c0",x"58",x"a6",x"d0"),
  2178 => (x"89",x"73",x"49",x"e0"),
  2179 => (x"28",x"71",x"48",x"74"),
  2180 => (x"c4",x"58",x"a6",x"d4"),
  2181 => (x"ba",x"ff",x"4a",x"66"),
  2182 => (x"66",x"c8",x"9a",x"6e"),
  2183 => (x"75",x"b9",x"ff",x"49"),
  2184 => (x"cc",x"48",x"72",x"99"),
  2185 => (x"c6",x"c3",x"b0",x"66"),
  2186 => (x"48",x"71",x"58",x"fe"),
  2187 => (x"c3",x"b0",x"66",x"d0"),
  2188 => (x"fb",x"58",x"c2",x"c7"),
  2189 => (x"8e",x"ec",x"87",x"c0"),
  2190 => (x"1e",x"87",x"f6",x"fc"),
  2191 => (x"c8",x"48",x"d0",x"ff"),
  2192 => (x"48",x"71",x"78",x"c9"),
  2193 => (x"78",x"08",x"d4",x"ff"),
  2194 => (x"71",x"1e",x"4f",x"26"),
  2195 => (x"87",x"eb",x"49",x"4a"),
  2196 => (x"c8",x"48",x"d0",x"ff"),
  2197 => (x"1e",x"4f",x"26",x"78"),
  2198 => (x"4b",x"71",x"1e",x"73"),
  2199 => (x"bf",x"ce",x"c7",x"c3"),
  2200 => (x"c2",x"87",x"c3",x"02"),
  2201 => (x"d0",x"ff",x"87",x"eb"),
  2202 => (x"78",x"c9",x"c8",x"48"),
  2203 => (x"e0",x"c0",x"49",x"73"),
  2204 => (x"48",x"d4",x"ff",x"b1"),
  2205 => (x"c7",x"c3",x"78",x"71"),
  2206 => (x"78",x"c0",x"48",x"c2"),
  2207 => (x"c5",x"02",x"66",x"c8"),
  2208 => (x"49",x"ff",x"c3",x"87"),
  2209 => (x"49",x"c0",x"87",x"c2"),
  2210 => (x"59",x"ca",x"c7",x"c3"),
  2211 => (x"c6",x"02",x"66",x"cc"),
  2212 => (x"d5",x"d5",x"c5",x"87"),
  2213 => (x"cf",x"87",x"c4",x"4a"),
  2214 => (x"c3",x"4a",x"ff",x"ff"),
  2215 => (x"c3",x"5a",x"ce",x"c7"),
  2216 => (x"c1",x"48",x"ce",x"c7"),
  2217 => (x"26",x"87",x"c4",x"78"),
  2218 => (x"26",x"4c",x"26",x"4d"),
  2219 => (x"0e",x"4f",x"26",x"4b"),
  2220 => (x"5d",x"5c",x"5b",x"5e"),
  2221 => (x"c3",x"4a",x"71",x"0e"),
  2222 => (x"4c",x"bf",x"ca",x"c7"),
  2223 => (x"cb",x"02",x"9a",x"72"),
  2224 => (x"91",x"c8",x"49",x"87"),
  2225 => (x"4b",x"cd",x"c9",x"c2"),
  2226 => (x"87",x"c4",x"83",x"71"),
  2227 => (x"4b",x"cd",x"cd",x"c2"),
  2228 => (x"49",x"13",x"4d",x"c0"),
  2229 => (x"c7",x"c3",x"99",x"74"),
  2230 => (x"ff",x"b9",x"bf",x"c6"),
  2231 => (x"78",x"71",x"48",x"d4"),
  2232 => (x"85",x"2c",x"b7",x"c1"),
  2233 => (x"04",x"ad",x"b7",x"c8"),
  2234 => (x"c7",x"c3",x"87",x"e8"),
  2235 => (x"c8",x"48",x"bf",x"c2"),
  2236 => (x"c6",x"c7",x"c3",x"80"),
  2237 => (x"87",x"ef",x"fe",x"58"),
  2238 => (x"71",x"1e",x"73",x"1e"),
  2239 => (x"9a",x"4a",x"13",x"4b"),
  2240 => (x"72",x"87",x"cb",x"02"),
  2241 => (x"87",x"e7",x"fe",x"49"),
  2242 => (x"05",x"9a",x"4a",x"13"),
  2243 => (x"da",x"fe",x"87",x"f5"),
  2244 => (x"c7",x"c3",x"1e",x"87"),
  2245 => (x"c3",x"49",x"bf",x"c2"),
  2246 => (x"c1",x"48",x"c2",x"c7"),
  2247 => (x"c0",x"c4",x"78",x"a1"),
  2248 => (x"db",x"03",x"a9",x"b7"),
  2249 => (x"48",x"d4",x"ff",x"87"),
  2250 => (x"bf",x"c6",x"c7",x"c3"),
  2251 => (x"c2",x"c7",x"c3",x"78"),
  2252 => (x"c7",x"c3",x"49",x"bf"),
  2253 => (x"a1",x"c1",x"48",x"c2"),
  2254 => (x"b7",x"c0",x"c4",x"78"),
  2255 => (x"87",x"e5",x"04",x"a9"),
  2256 => (x"c8",x"48",x"d0",x"ff"),
  2257 => (x"ce",x"c7",x"c3",x"78"),
  2258 => (x"26",x"78",x"c0",x"48"),
  2259 => (x"00",x"00",x"00",x"4f"),
  2260 => (x"00",x"00",x"00",x"00"),
  2261 => (x"00",x"00",x"00",x"00"),
  2262 => (x"00",x"00",x"5f",x"5f"),
  2263 => (x"03",x"03",x"00",x"00"),
  2264 => (x"00",x"03",x"03",x"00"),
  2265 => (x"7f",x"7f",x"14",x"00"),
  2266 => (x"14",x"7f",x"7f",x"14"),
  2267 => (x"2e",x"24",x"00",x"00"),
  2268 => (x"12",x"3a",x"6b",x"6b"),
  2269 => (x"36",x"6a",x"4c",x"00"),
  2270 => (x"32",x"56",x"6c",x"18"),
  2271 => (x"4f",x"7e",x"30",x"00"),
  2272 => (x"68",x"3a",x"77",x"59"),
  2273 => (x"04",x"00",x"00",x"40"),
  2274 => (x"00",x"00",x"03",x"07"),
  2275 => (x"1c",x"00",x"00",x"00"),
  2276 => (x"00",x"41",x"63",x"3e"),
  2277 => (x"41",x"00",x"00",x"00"),
  2278 => (x"00",x"1c",x"3e",x"63"),
  2279 => (x"3e",x"2a",x"08",x"00"),
  2280 => (x"2a",x"3e",x"1c",x"1c"),
  2281 => (x"08",x"08",x"00",x"08"),
  2282 => (x"08",x"08",x"3e",x"3e"),
  2283 => (x"80",x"00",x"00",x"00"),
  2284 => (x"00",x"00",x"60",x"e0"),
  2285 => (x"08",x"08",x"00",x"00"),
  2286 => (x"08",x"08",x"08",x"08"),
  2287 => (x"00",x"00",x"00",x"00"),
  2288 => (x"00",x"00",x"60",x"60"),
  2289 => (x"30",x"60",x"40",x"00"),
  2290 => (x"03",x"06",x"0c",x"18"),
  2291 => (x"7f",x"3e",x"00",x"01"),
  2292 => (x"3e",x"7f",x"4d",x"59"),
  2293 => (x"06",x"04",x"00",x"00"),
  2294 => (x"00",x"00",x"7f",x"7f"),
  2295 => (x"63",x"42",x"00",x"00"),
  2296 => (x"46",x"4f",x"59",x"71"),
  2297 => (x"63",x"22",x"00",x"00"),
  2298 => (x"36",x"7f",x"49",x"49"),
  2299 => (x"16",x"1c",x"18",x"00"),
  2300 => (x"10",x"7f",x"7f",x"13"),
  2301 => (x"67",x"27",x"00",x"00"),
  2302 => (x"39",x"7d",x"45",x"45"),
  2303 => (x"7e",x"3c",x"00",x"00"),
  2304 => (x"30",x"79",x"49",x"4b"),
  2305 => (x"01",x"01",x"00",x"00"),
  2306 => (x"07",x"0f",x"79",x"71"),
  2307 => (x"7f",x"36",x"00",x"00"),
  2308 => (x"36",x"7f",x"49",x"49"),
  2309 => (x"4f",x"06",x"00",x"00"),
  2310 => (x"1e",x"3f",x"69",x"49"),
  2311 => (x"00",x"00",x"00",x"00"),
  2312 => (x"00",x"00",x"66",x"66"),
  2313 => (x"80",x"00",x"00",x"00"),
  2314 => (x"00",x"00",x"66",x"e6"),
  2315 => (x"08",x"08",x"00",x"00"),
  2316 => (x"22",x"22",x"14",x"14"),
  2317 => (x"14",x"14",x"00",x"00"),
  2318 => (x"14",x"14",x"14",x"14"),
  2319 => (x"22",x"22",x"00",x"00"),
  2320 => (x"08",x"08",x"14",x"14"),
  2321 => (x"03",x"02",x"00",x"00"),
  2322 => (x"06",x"0f",x"59",x"51"),
  2323 => (x"41",x"7f",x"3e",x"00"),
  2324 => (x"1e",x"1f",x"55",x"5d"),
  2325 => (x"7f",x"7e",x"00",x"00"),
  2326 => (x"7e",x"7f",x"09",x"09"),
  2327 => (x"7f",x"7f",x"00",x"00"),
  2328 => (x"36",x"7f",x"49",x"49"),
  2329 => (x"3e",x"1c",x"00",x"00"),
  2330 => (x"41",x"41",x"41",x"63"),
  2331 => (x"7f",x"7f",x"00",x"00"),
  2332 => (x"1c",x"3e",x"63",x"41"),
  2333 => (x"7f",x"7f",x"00",x"00"),
  2334 => (x"41",x"41",x"49",x"49"),
  2335 => (x"7f",x"7f",x"00",x"00"),
  2336 => (x"01",x"01",x"09",x"09"),
  2337 => (x"7f",x"3e",x"00",x"00"),
  2338 => (x"7a",x"7b",x"49",x"41"),
  2339 => (x"7f",x"7f",x"00",x"00"),
  2340 => (x"7f",x"7f",x"08",x"08"),
  2341 => (x"41",x"00",x"00",x"00"),
  2342 => (x"00",x"41",x"7f",x"7f"),
  2343 => (x"60",x"20",x"00",x"00"),
  2344 => (x"3f",x"7f",x"40",x"40"),
  2345 => (x"08",x"7f",x"7f",x"00"),
  2346 => (x"41",x"63",x"36",x"1c"),
  2347 => (x"7f",x"7f",x"00",x"00"),
  2348 => (x"40",x"40",x"40",x"40"),
  2349 => (x"06",x"7f",x"7f",x"00"),
  2350 => (x"7f",x"7f",x"06",x"0c"),
  2351 => (x"06",x"7f",x"7f",x"00"),
  2352 => (x"7f",x"7f",x"18",x"0c"),
  2353 => (x"7f",x"3e",x"00",x"00"),
  2354 => (x"3e",x"7f",x"41",x"41"),
  2355 => (x"7f",x"7f",x"00",x"00"),
  2356 => (x"06",x"0f",x"09",x"09"),
  2357 => (x"41",x"7f",x"3e",x"00"),
  2358 => (x"40",x"7e",x"7f",x"61"),
  2359 => (x"7f",x"7f",x"00",x"00"),
  2360 => (x"66",x"7f",x"19",x"09"),
  2361 => (x"6f",x"26",x"00",x"00"),
  2362 => (x"32",x"7b",x"59",x"4d"),
  2363 => (x"01",x"01",x"00",x"00"),
  2364 => (x"01",x"01",x"7f",x"7f"),
  2365 => (x"7f",x"3f",x"00",x"00"),
  2366 => (x"3f",x"7f",x"40",x"40"),
  2367 => (x"3f",x"0f",x"00",x"00"),
  2368 => (x"0f",x"3f",x"70",x"70"),
  2369 => (x"30",x"7f",x"7f",x"00"),
  2370 => (x"7f",x"7f",x"30",x"18"),
  2371 => (x"36",x"63",x"41",x"00"),
  2372 => (x"63",x"36",x"1c",x"1c"),
  2373 => (x"06",x"03",x"01",x"41"),
  2374 => (x"03",x"06",x"7c",x"7c"),
  2375 => (x"59",x"71",x"61",x"01"),
  2376 => (x"41",x"43",x"47",x"4d"),
  2377 => (x"7f",x"00",x"00",x"00"),
  2378 => (x"00",x"41",x"41",x"7f"),
  2379 => (x"06",x"03",x"01",x"00"),
  2380 => (x"60",x"30",x"18",x"0c"),
  2381 => (x"41",x"00",x"00",x"40"),
  2382 => (x"00",x"7f",x"7f",x"41"),
  2383 => (x"06",x"0c",x"08",x"00"),
  2384 => (x"08",x"0c",x"06",x"03"),
  2385 => (x"80",x"80",x"80",x"00"),
  2386 => (x"80",x"80",x"80",x"80"),
  2387 => (x"00",x"00",x"00",x"00"),
  2388 => (x"00",x"04",x"07",x"03"),
  2389 => (x"74",x"20",x"00",x"00"),
  2390 => (x"78",x"7c",x"54",x"54"),
  2391 => (x"7f",x"7f",x"00",x"00"),
  2392 => (x"38",x"7c",x"44",x"44"),
  2393 => (x"7c",x"38",x"00",x"00"),
  2394 => (x"00",x"44",x"44",x"44"),
  2395 => (x"7c",x"38",x"00",x"00"),
  2396 => (x"7f",x"7f",x"44",x"44"),
  2397 => (x"7c",x"38",x"00",x"00"),
  2398 => (x"18",x"5c",x"54",x"54"),
  2399 => (x"7e",x"04",x"00",x"00"),
  2400 => (x"00",x"05",x"05",x"7f"),
  2401 => (x"bc",x"18",x"00",x"00"),
  2402 => (x"7c",x"fc",x"a4",x"a4"),
  2403 => (x"7f",x"7f",x"00",x"00"),
  2404 => (x"78",x"7c",x"04",x"04"),
  2405 => (x"00",x"00",x"00",x"00"),
  2406 => (x"00",x"40",x"7d",x"3d"),
  2407 => (x"80",x"80",x"00",x"00"),
  2408 => (x"00",x"7d",x"fd",x"80"),
  2409 => (x"7f",x"7f",x"00",x"00"),
  2410 => (x"44",x"6c",x"38",x"10"),
  2411 => (x"00",x"00",x"00",x"00"),
  2412 => (x"00",x"40",x"7f",x"3f"),
  2413 => (x"0c",x"7c",x"7c",x"00"),
  2414 => (x"78",x"7c",x"0c",x"18"),
  2415 => (x"7c",x"7c",x"00",x"00"),
  2416 => (x"78",x"7c",x"04",x"04"),
  2417 => (x"7c",x"38",x"00",x"00"),
  2418 => (x"38",x"7c",x"44",x"44"),
  2419 => (x"fc",x"fc",x"00",x"00"),
  2420 => (x"18",x"3c",x"24",x"24"),
  2421 => (x"3c",x"18",x"00",x"00"),
  2422 => (x"fc",x"fc",x"24",x"24"),
  2423 => (x"7c",x"7c",x"00",x"00"),
  2424 => (x"08",x"0c",x"04",x"04"),
  2425 => (x"5c",x"48",x"00",x"00"),
  2426 => (x"20",x"74",x"54",x"54"),
  2427 => (x"3f",x"04",x"00",x"00"),
  2428 => (x"00",x"44",x"44",x"7f"),
  2429 => (x"7c",x"3c",x"00",x"00"),
  2430 => (x"7c",x"7c",x"40",x"40"),
  2431 => (x"3c",x"1c",x"00",x"00"),
  2432 => (x"1c",x"3c",x"60",x"60"),
  2433 => (x"60",x"7c",x"3c",x"00"),
  2434 => (x"3c",x"7c",x"60",x"30"),
  2435 => (x"38",x"6c",x"44",x"00"),
  2436 => (x"44",x"6c",x"38",x"10"),
  2437 => (x"bc",x"1c",x"00",x"00"),
  2438 => (x"1c",x"3c",x"60",x"e0"),
  2439 => (x"64",x"44",x"00",x"00"),
  2440 => (x"44",x"4c",x"5c",x"74"),
  2441 => (x"08",x"08",x"00",x"00"),
  2442 => (x"41",x"41",x"77",x"3e"),
  2443 => (x"00",x"00",x"00",x"00"),
  2444 => (x"00",x"00",x"7f",x"7f"),
  2445 => (x"41",x"41",x"00",x"00"),
  2446 => (x"08",x"08",x"3e",x"77"),
  2447 => (x"01",x"01",x"02",x"00"),
  2448 => (x"01",x"02",x"02",x"03"),
  2449 => (x"7f",x"7f",x"7f",x"00"),
  2450 => (x"7f",x"7f",x"7f",x"7f"),
  2451 => (x"1c",x"08",x"08",x"00"),
  2452 => (x"7f",x"3e",x"3e",x"1c"),
  2453 => (x"3e",x"7f",x"7f",x"7f"),
  2454 => (x"08",x"1c",x"1c",x"3e"),
  2455 => (x"18",x"10",x"00",x"08"),
  2456 => (x"10",x"18",x"7c",x"7c"),
  2457 => (x"30",x"10",x"00",x"00"),
  2458 => (x"10",x"30",x"7c",x"7c"),
  2459 => (x"60",x"30",x"10",x"00"),
  2460 => (x"06",x"1e",x"78",x"60"),
  2461 => (x"3c",x"66",x"42",x"00"),
  2462 => (x"42",x"66",x"3c",x"18"),
  2463 => (x"6a",x"38",x"78",x"00"),
  2464 => (x"38",x"6c",x"c6",x"c2"),
  2465 => (x"00",x"00",x"60",x"00"),
  2466 => (x"60",x"00",x"00",x"60"),
  2467 => (x"5b",x"5e",x"0e",x"00"),
  2468 => (x"1e",x"0e",x"5d",x"5c"),
  2469 => (x"c7",x"c3",x"4c",x"71"),
  2470 => (x"c0",x"4d",x"bf",x"df"),
  2471 => (x"74",x"1e",x"c0",x"4b"),
  2472 => (x"87",x"c7",x"02",x"ab"),
  2473 => (x"c0",x"48",x"a6",x"c4"),
  2474 => (x"c4",x"87",x"c5",x"78"),
  2475 => (x"78",x"c1",x"48",x"a6"),
  2476 => (x"73",x"1e",x"66",x"c4"),
  2477 => (x"87",x"df",x"ee",x"49"),
  2478 => (x"e0",x"c0",x"86",x"c8"),
  2479 => (x"87",x"ef",x"ef",x"49"),
  2480 => (x"6a",x"4a",x"a5",x"c4"),
  2481 => (x"87",x"f0",x"f0",x"49"),
  2482 => (x"cb",x"87",x"c6",x"f1"),
  2483 => (x"c8",x"83",x"c1",x"85"),
  2484 => (x"ff",x"04",x"ab",x"b7"),
  2485 => (x"26",x"26",x"87",x"c7"),
  2486 => (x"26",x"4c",x"26",x"4d"),
  2487 => (x"1e",x"4f",x"26",x"4b"),
  2488 => (x"c7",x"c3",x"4a",x"71"),
  2489 => (x"c7",x"c3",x"5a",x"e3"),
  2490 => (x"78",x"c7",x"48",x"e3"),
  2491 => (x"87",x"dd",x"fe",x"49"),
  2492 => (x"73",x"1e",x"4f",x"26"),
  2493 => (x"c0",x"4a",x"71",x"1e"),
  2494 => (x"d3",x"03",x"aa",x"b7"),
  2495 => (x"d1",x"e9",x"c2",x"87"),
  2496 => (x"87",x"c4",x"05",x"bf"),
  2497 => (x"87",x"c2",x"4b",x"c1"),
  2498 => (x"e9",x"c2",x"4b",x"c0"),
  2499 => (x"87",x"c4",x"5b",x"d5"),
  2500 => (x"5a",x"d5",x"e9",x"c2"),
  2501 => (x"bf",x"d1",x"e9",x"c2"),
  2502 => (x"c1",x"9a",x"c1",x"4a"),
  2503 => (x"ec",x"49",x"a2",x"c0"),
  2504 => (x"48",x"fc",x"87",x"e8"),
  2505 => (x"bf",x"d1",x"e9",x"c2"),
  2506 => (x"87",x"ef",x"fe",x"78"),
  2507 => (x"c4",x"4a",x"71",x"1e"),
  2508 => (x"49",x"72",x"1e",x"66"),
  2509 => (x"26",x"87",x"e2",x"e6"),
  2510 => (x"c2",x"1e",x"4f",x"26"),
  2511 => (x"49",x"bf",x"d1",x"e9"),
  2512 => (x"87",x"f2",x"da",x"ff"),
  2513 => (x"48",x"d7",x"c7",x"c3"),
  2514 => (x"c3",x"78",x"bf",x"e8"),
  2515 => (x"ec",x"48",x"d3",x"c7"),
  2516 => (x"c7",x"c3",x"78",x"bf"),
  2517 => (x"49",x"4a",x"bf",x"d7"),
  2518 => (x"c8",x"99",x"ff",x"c3"),
  2519 => (x"48",x"72",x"2a",x"b7"),
  2520 => (x"c7",x"c3",x"b0",x"71"),
  2521 => (x"4f",x"26",x"58",x"df"),
  2522 => (x"5c",x"5b",x"5e",x"0e"),
  2523 => (x"4b",x"71",x"0e",x"5d"),
  2524 => (x"c3",x"87",x"c7",x"ff"),
  2525 => (x"c0",x"48",x"d2",x"c7"),
  2526 => (x"ff",x"49",x"73",x"50"),
  2527 => (x"70",x"87",x"d7",x"da"),
  2528 => (x"9c",x"c2",x"4c",x"49"),
  2529 => (x"cb",x"49",x"ee",x"cb"),
  2530 => (x"49",x"70",x"87",x"cf"),
  2531 => (x"d2",x"c7",x"c3",x"4d"),
  2532 => (x"c1",x"05",x"bf",x"97"),
  2533 => (x"66",x"d0",x"87",x"e4"),
  2534 => (x"db",x"c7",x"c3",x"49"),
  2535 => (x"d7",x"05",x"99",x"bf"),
  2536 => (x"49",x"66",x"d4",x"87"),
  2537 => (x"bf",x"d3",x"c7",x"c3"),
  2538 => (x"87",x"cc",x"05",x"99"),
  2539 => (x"d9",x"ff",x"49",x"73"),
  2540 => (x"98",x"70",x"87",x"e4"),
  2541 => (x"87",x"c2",x"c1",x"02"),
  2542 => (x"fd",x"fd",x"4c",x"c1"),
  2543 => (x"ca",x"49",x"75",x"87"),
  2544 => (x"98",x"70",x"87",x"e3"),
  2545 => (x"c3",x"87",x"c6",x"02"),
  2546 => (x"c1",x"48",x"d2",x"c7"),
  2547 => (x"d2",x"c7",x"c3",x"50"),
  2548 => (x"c0",x"05",x"bf",x"97"),
  2549 => (x"c7",x"c3",x"87",x"e4"),
  2550 => (x"d0",x"49",x"bf",x"db"),
  2551 => (x"ff",x"05",x"99",x"66"),
  2552 => (x"c7",x"c3",x"87",x"d6"),
  2553 => (x"d4",x"49",x"bf",x"d3"),
  2554 => (x"ff",x"05",x"99",x"66"),
  2555 => (x"49",x"73",x"87",x"ca"),
  2556 => (x"87",x"e2",x"d8",x"ff"),
  2557 => (x"fe",x"05",x"98",x"70"),
  2558 => (x"48",x"74",x"87",x"fe"),
  2559 => (x"0e",x"87",x"d8",x"fb"),
  2560 => (x"5d",x"5c",x"5b",x"5e"),
  2561 => (x"c0",x"86",x"f4",x"0e"),
  2562 => (x"bf",x"ec",x"4c",x"4d"),
  2563 => (x"48",x"a6",x"c4",x"7e"),
  2564 => (x"bf",x"df",x"c7",x"c3"),
  2565 => (x"c0",x"1e",x"c1",x"78"),
  2566 => (x"fd",x"49",x"c7",x"1e"),
  2567 => (x"86",x"c8",x"87",x"ca"),
  2568 => (x"ce",x"02",x"98",x"70"),
  2569 => (x"fb",x"49",x"ff",x"87"),
  2570 => (x"da",x"c1",x"87",x"c8"),
  2571 => (x"e5",x"d7",x"ff",x"49"),
  2572 => (x"c3",x"4d",x"c1",x"87"),
  2573 => (x"bf",x"97",x"d2",x"c7"),
  2574 => (x"d0",x"87",x"c3",x"02"),
  2575 => (x"c7",x"c3",x"87",x"c5"),
  2576 => (x"c2",x"4b",x"bf",x"d7"),
  2577 => (x"05",x"bf",x"d1",x"e9"),
  2578 => (x"c3",x"87",x"eb",x"c0"),
  2579 => (x"d7",x"ff",x"49",x"fd"),
  2580 => (x"fa",x"c3",x"87",x"c4"),
  2581 => (x"fd",x"d6",x"ff",x"49"),
  2582 => (x"c3",x"49",x"73",x"87"),
  2583 => (x"1e",x"71",x"99",x"ff"),
  2584 => (x"c7",x"fb",x"49",x"c0"),
  2585 => (x"c8",x"49",x"73",x"87"),
  2586 => (x"1e",x"71",x"29",x"b7"),
  2587 => (x"fb",x"fa",x"49",x"c1"),
  2588 => (x"c6",x"86",x"c8",x"87"),
  2589 => (x"c7",x"c3",x"87",x"c1"),
  2590 => (x"9b",x"4b",x"bf",x"db"),
  2591 => (x"c2",x"87",x"dd",x"02"),
  2592 => (x"49",x"bf",x"cd",x"e9"),
  2593 => (x"70",x"87",x"de",x"c7"),
  2594 => (x"87",x"c4",x"05",x"98"),
  2595 => (x"87",x"d2",x"4b",x"c0"),
  2596 => (x"c7",x"49",x"e0",x"c2"),
  2597 => (x"e9",x"c2",x"87",x"c3"),
  2598 => (x"87",x"c6",x"58",x"d1"),
  2599 => (x"48",x"cd",x"e9",x"c2"),
  2600 => (x"49",x"73",x"78",x"c0"),
  2601 => (x"ce",x"05",x"99",x"c2"),
  2602 => (x"49",x"eb",x"c3",x"87"),
  2603 => (x"87",x"e6",x"d5",x"ff"),
  2604 => (x"99",x"c2",x"49",x"70"),
  2605 => (x"fb",x"87",x"c2",x"02"),
  2606 => (x"c1",x"49",x"73",x"4c"),
  2607 => (x"87",x"ce",x"05",x"99"),
  2608 => (x"ff",x"49",x"f4",x"c3"),
  2609 => (x"70",x"87",x"cf",x"d5"),
  2610 => (x"02",x"99",x"c2",x"49"),
  2611 => (x"4c",x"fa",x"87",x"c2"),
  2612 => (x"99",x"c8",x"49",x"73"),
  2613 => (x"c3",x"87",x"ce",x"05"),
  2614 => (x"d4",x"ff",x"49",x"f5"),
  2615 => (x"49",x"70",x"87",x"f8"),
  2616 => (x"d5",x"02",x"99",x"c2"),
  2617 => (x"e3",x"c7",x"c3",x"87"),
  2618 => (x"87",x"ca",x"02",x"bf"),
  2619 => (x"c3",x"88",x"c1",x"48"),
  2620 => (x"c0",x"58",x"e7",x"c7"),
  2621 => (x"4c",x"ff",x"87",x"c2"),
  2622 => (x"49",x"73",x"4d",x"c1"),
  2623 => (x"ce",x"05",x"99",x"c4"),
  2624 => (x"49",x"f2",x"c3",x"87"),
  2625 => (x"87",x"ce",x"d4",x"ff"),
  2626 => (x"99",x"c2",x"49",x"70"),
  2627 => (x"c3",x"87",x"dc",x"02"),
  2628 => (x"7e",x"bf",x"e3",x"c7"),
  2629 => (x"a8",x"b7",x"c7",x"48"),
  2630 => (x"87",x"cb",x"c0",x"03"),
  2631 => (x"80",x"c1",x"48",x"6e"),
  2632 => (x"58",x"e7",x"c7",x"c3"),
  2633 => (x"fe",x"87",x"c2",x"c0"),
  2634 => (x"c3",x"4d",x"c1",x"4c"),
  2635 => (x"d3",x"ff",x"49",x"fd"),
  2636 => (x"49",x"70",x"87",x"e4"),
  2637 => (x"c0",x"02",x"99",x"c2"),
  2638 => (x"c7",x"c3",x"87",x"d5"),
  2639 => (x"c0",x"02",x"bf",x"e3"),
  2640 => (x"c7",x"c3",x"87",x"c9"),
  2641 => (x"78",x"c0",x"48",x"e3"),
  2642 => (x"fd",x"87",x"c2",x"c0"),
  2643 => (x"c3",x"4d",x"c1",x"4c"),
  2644 => (x"d3",x"ff",x"49",x"fa"),
  2645 => (x"49",x"70",x"87",x"c0"),
  2646 => (x"c0",x"02",x"99",x"c2"),
  2647 => (x"c7",x"c3",x"87",x"d9"),
  2648 => (x"c7",x"48",x"bf",x"e3"),
  2649 => (x"c0",x"03",x"a8",x"b7"),
  2650 => (x"c7",x"c3",x"87",x"c9"),
  2651 => (x"78",x"c7",x"48",x"e3"),
  2652 => (x"fc",x"87",x"c2",x"c0"),
  2653 => (x"c0",x"4d",x"c1",x"4c"),
  2654 => (x"c0",x"03",x"ac",x"b7"),
  2655 => (x"66",x"c4",x"87",x"d1"),
  2656 => (x"82",x"d8",x"c1",x"4a"),
  2657 => (x"c6",x"c0",x"02",x"6a"),
  2658 => (x"74",x"4b",x"6a",x"87"),
  2659 => (x"c0",x"0f",x"73",x"49"),
  2660 => (x"1e",x"f0",x"c3",x"1e"),
  2661 => (x"f7",x"49",x"da",x"c1"),
  2662 => (x"86",x"c8",x"87",x"ce"),
  2663 => (x"c0",x"02",x"98",x"70"),
  2664 => (x"a6",x"c8",x"87",x"e2"),
  2665 => (x"e3",x"c7",x"c3",x"48"),
  2666 => (x"66",x"c8",x"78",x"bf"),
  2667 => (x"c4",x"91",x"cb",x"49"),
  2668 => (x"80",x"71",x"48",x"66"),
  2669 => (x"bf",x"6e",x"7e",x"70"),
  2670 => (x"87",x"c8",x"c0",x"02"),
  2671 => (x"c8",x"4b",x"bf",x"6e"),
  2672 => (x"0f",x"73",x"49",x"66"),
  2673 => (x"c0",x"02",x"9d",x"75"),
  2674 => (x"c7",x"c3",x"87",x"c8"),
  2675 => (x"f2",x"49",x"bf",x"e3"),
  2676 => (x"e9",x"c2",x"87",x"fb"),
  2677 => (x"c0",x"02",x"bf",x"d5"),
  2678 => (x"c2",x"49",x"87",x"dd"),
  2679 => (x"98",x"70",x"87",x"c7"),
  2680 => (x"87",x"d3",x"c0",x"02"),
  2681 => (x"bf",x"e3",x"c7",x"c3"),
  2682 => (x"87",x"e1",x"f2",x"49"),
  2683 => (x"c1",x"f4",x"49",x"c0"),
  2684 => (x"d5",x"e9",x"c2",x"87"),
  2685 => (x"f4",x"78",x"c0",x"48"),
  2686 => (x"87",x"db",x"f3",x"8e"),
  2687 => (x"5c",x"5b",x"5e",x"0e"),
  2688 => (x"71",x"1e",x"0e",x"5d"),
  2689 => (x"df",x"c7",x"c3",x"4c"),
  2690 => (x"cd",x"c1",x"49",x"bf"),
  2691 => (x"d1",x"c1",x"4d",x"a1"),
  2692 => (x"74",x"7e",x"69",x"81"),
  2693 => (x"87",x"cf",x"02",x"9c"),
  2694 => (x"74",x"4b",x"a5",x"c4"),
  2695 => (x"df",x"c7",x"c3",x"7b"),
  2696 => (x"fa",x"f2",x"49",x"bf"),
  2697 => (x"74",x"7b",x"6e",x"87"),
  2698 => (x"87",x"c4",x"05",x"9c"),
  2699 => (x"87",x"c2",x"4b",x"c0"),
  2700 => (x"49",x"73",x"4b",x"c1"),
  2701 => (x"d4",x"87",x"fb",x"f2"),
  2702 => (x"87",x"c7",x"02",x"66"),
  2703 => (x"70",x"87",x"da",x"49"),
  2704 => (x"c0",x"87",x"c2",x"4a"),
  2705 => (x"d9",x"e9",x"c2",x"4a"),
  2706 => (x"ca",x"f2",x"26",x"5a"),
  2707 => (x"00",x"00",x"00",x"87"),
  2708 => (x"00",x"00",x"00",x"00"),
  2709 => (x"00",x"00",x"00",x"00"),
  2710 => (x"4a",x"71",x"1e",x"00"),
  2711 => (x"49",x"bf",x"c8",x"ff"),
  2712 => (x"26",x"48",x"a1",x"72"),
  2713 => (x"c8",x"ff",x"1e",x"4f"),
  2714 => (x"c0",x"fe",x"89",x"bf"),
  2715 => (x"c0",x"c0",x"c0",x"c0"),
  2716 => (x"87",x"c4",x"01",x"a9"),
  2717 => (x"87",x"c2",x"4a",x"c0"),
  2718 => (x"48",x"72",x"4a",x"c1"),
  2719 => (x"5e",x"0e",x"4f",x"26"),
  2720 => (x"0e",x"5d",x"5c",x"5b"),
  2721 => (x"d4",x"ff",x"4b",x"71"),
  2722 => (x"48",x"66",x"d0",x"4c"),
  2723 => (x"49",x"d6",x"78",x"c0"),
  2724 => (x"87",x"cb",x"d8",x"ff"),
  2725 => (x"6c",x"7c",x"ff",x"c3"),
  2726 => (x"99",x"ff",x"c3",x"49"),
  2727 => (x"c3",x"49",x"4d",x"71"),
  2728 => (x"e0",x"c1",x"99",x"f0"),
  2729 => (x"87",x"cb",x"05",x"a9"),
  2730 => (x"6c",x"7c",x"ff",x"c3"),
  2731 => (x"d0",x"98",x"c3",x"48"),
  2732 => (x"c3",x"78",x"08",x"66"),
  2733 => (x"4a",x"6c",x"7c",x"ff"),
  2734 => (x"c3",x"31",x"c8",x"49"),
  2735 => (x"4a",x"6c",x"7c",x"ff"),
  2736 => (x"49",x"72",x"b2",x"71"),
  2737 => (x"ff",x"c3",x"31",x"c8"),
  2738 => (x"71",x"4a",x"6c",x"7c"),
  2739 => (x"c8",x"49",x"72",x"b2"),
  2740 => (x"7c",x"ff",x"c3",x"31"),
  2741 => (x"b2",x"71",x"4a",x"6c"),
  2742 => (x"c0",x"48",x"d0",x"ff"),
  2743 => (x"9b",x"73",x"78",x"e0"),
  2744 => (x"72",x"87",x"c2",x"02"),
  2745 => (x"26",x"48",x"75",x"7b"),
  2746 => (x"26",x"4c",x"26",x"4d"),
  2747 => (x"1e",x"4f",x"26",x"4b"),
  2748 => (x"5e",x"0e",x"4f",x"26"),
  2749 => (x"f8",x"0e",x"5c",x"5b"),
  2750 => (x"c8",x"1e",x"76",x"86"),
  2751 => (x"fd",x"fd",x"49",x"a6"),
  2752 => (x"70",x"86",x"c4",x"87"),
  2753 => (x"c2",x"48",x"6e",x"4b"),
  2754 => (x"f0",x"c2",x"03",x"a8"),
  2755 => (x"c3",x"4a",x"73",x"87"),
  2756 => (x"d0",x"c1",x"9a",x"f0"),
  2757 => (x"87",x"c7",x"02",x"aa"),
  2758 => (x"05",x"aa",x"e0",x"c1"),
  2759 => (x"73",x"87",x"de",x"c2"),
  2760 => (x"02",x"99",x"c8",x"49"),
  2761 => (x"c6",x"ff",x"87",x"c3"),
  2762 => (x"c3",x"4c",x"73",x"87"),
  2763 => (x"05",x"ac",x"c2",x"9c"),
  2764 => (x"c4",x"87",x"c2",x"c1"),
  2765 => (x"31",x"c9",x"49",x"66"),
  2766 => (x"66",x"c4",x"1e",x"71"),
  2767 => (x"c3",x"92",x"d4",x"4a"),
  2768 => (x"72",x"49",x"e7",x"c7"),
  2769 => (x"d7",x"fa",x"fd",x"81"),
  2770 => (x"ff",x"49",x"d8",x"87"),
  2771 => (x"c8",x"87",x"d0",x"d5"),
  2772 => (x"f5",x"c2",x"1e",x"c0"),
  2773 => (x"d6",x"fd",x"49",x"de"),
  2774 => (x"d0",x"ff",x"87",x"d2"),
  2775 => (x"78",x"e0",x"c0",x"48"),
  2776 => (x"1e",x"de",x"f5",x"c2"),
  2777 => (x"d4",x"4a",x"66",x"cc"),
  2778 => (x"e7",x"c7",x"c3",x"92"),
  2779 => (x"fd",x"81",x"72",x"49"),
  2780 => (x"cc",x"87",x"de",x"f8"),
  2781 => (x"05",x"ac",x"c1",x"86"),
  2782 => (x"c4",x"87",x"c2",x"c1"),
  2783 => (x"31",x"c9",x"49",x"66"),
  2784 => (x"66",x"c4",x"1e",x"71"),
  2785 => (x"c3",x"92",x"d4",x"4a"),
  2786 => (x"72",x"49",x"e7",x"c7"),
  2787 => (x"cf",x"f9",x"fd",x"81"),
  2788 => (x"de",x"f5",x"c2",x"87"),
  2789 => (x"4a",x"66",x"c8",x"1e"),
  2790 => (x"c7",x"c3",x"92",x"d4"),
  2791 => (x"81",x"72",x"49",x"e7"),
  2792 => (x"87",x"de",x"f6",x"fd"),
  2793 => (x"d3",x"ff",x"49",x"d7"),
  2794 => (x"c0",x"c8",x"87",x"f5"),
  2795 => (x"de",x"f5",x"c2",x"1e"),
  2796 => (x"d0",x"d4",x"fd",x"49"),
  2797 => (x"ff",x"86",x"cc",x"87"),
  2798 => (x"e0",x"c0",x"48",x"d0"),
  2799 => (x"fc",x"8e",x"f8",x"78"),
  2800 => (x"5e",x"0e",x"87",x"e7"),
  2801 => (x"0e",x"5d",x"5c",x"5b"),
  2802 => (x"ff",x"4d",x"71",x"1e"),
  2803 => (x"66",x"d4",x"4c",x"d4"),
  2804 => (x"b7",x"c3",x"48",x"7e"),
  2805 => (x"87",x"c5",x"06",x"a8"),
  2806 => (x"e2",x"c1",x"48",x"c0"),
  2807 => (x"fe",x"49",x"75",x"87"),
  2808 => (x"75",x"87",x"e3",x"c7"),
  2809 => (x"4b",x"66",x"c4",x"1e"),
  2810 => (x"c7",x"c3",x"93",x"d4"),
  2811 => (x"49",x"73",x"83",x"e7"),
  2812 => (x"87",x"f9",x"f1",x"fd"),
  2813 => (x"4b",x"6b",x"83",x"c8"),
  2814 => (x"c8",x"48",x"d0",x"ff"),
  2815 => (x"7c",x"dd",x"78",x"e1"),
  2816 => (x"ff",x"c3",x"49",x"73"),
  2817 => (x"73",x"7c",x"71",x"99"),
  2818 => (x"29",x"b7",x"c8",x"49"),
  2819 => (x"71",x"99",x"ff",x"c3"),
  2820 => (x"d0",x"49",x"73",x"7c"),
  2821 => (x"ff",x"c3",x"29",x"b7"),
  2822 => (x"73",x"7c",x"71",x"99"),
  2823 => (x"29",x"b7",x"d8",x"49"),
  2824 => (x"7c",x"c0",x"7c",x"71"),
  2825 => (x"7c",x"7c",x"7c",x"7c"),
  2826 => (x"7c",x"7c",x"7c",x"7c"),
  2827 => (x"c0",x"7c",x"7c",x"7c"),
  2828 => (x"66",x"c4",x"78",x"e0"),
  2829 => (x"ff",x"49",x"dc",x"1e"),
  2830 => (x"c8",x"87",x"c9",x"d2"),
  2831 => (x"26",x"48",x"73",x"86"),
  2832 => (x"1e",x"87",x"e4",x"fa"),
  2833 => (x"bf",x"f4",x"f4",x"c2"),
  2834 => (x"c2",x"b9",x"c1",x"49"),
  2835 => (x"ff",x"59",x"f8",x"f4"),
  2836 => (x"ff",x"c3",x"48",x"d4"),
  2837 => (x"48",x"d0",x"ff",x"78"),
  2838 => (x"ff",x"78",x"e1",x"c8"),
  2839 => (x"78",x"c1",x"48",x"d4"),
  2840 => (x"78",x"71",x"31",x"c4"),
  2841 => (x"c0",x"48",x"d0",x"ff"),
  2842 => (x"4f",x"26",x"78",x"e0"),
  2843 => (x"c5",x"f2",x"c2",x"1e"),
  2844 => (x"d4",x"c2",x"c3",x"1e"),
  2845 => (x"f4",x"ef",x"fd",x"49"),
  2846 => (x"70",x"86",x"c4",x"87"),
  2847 => (x"87",x"c3",x"02",x"98"),
  2848 => (x"26",x"87",x"c0",x"ff"),
  2849 => (x"4b",x"35",x"31",x"4f"),
  2850 => (x"20",x"20",x"5a",x"48"),
  2851 => (x"47",x"46",x"43",x"20"),
  2852 => (x"4a",x"71",x"1e",x"00"),
  2853 => (x"c3",x"49",x"a2",x"c4"),
  2854 => (x"6a",x"48",x"fa",x"c6"),
  2855 => (x"c1",x"49",x"69",x"78"),
  2856 => (x"f8",x"f4",x"c2",x"b9"),
  2857 => (x"87",x"db",x"fe",x"59"),
  2858 => (x"87",x"ca",x"d1",x"ff"),
  2859 => (x"4f",x"26",x"48",x"c1"),
  2860 => (x"c4",x"4a",x"71",x"1e"),
  2861 => (x"c6",x"c3",x"49",x"a2"),
  2862 => (x"c2",x"7a",x"bf",x"fa"),
  2863 => (x"79",x"bf",x"f4",x"f4"),
  2864 => (x"71",x"1e",x"4f",x"26"),
  2865 => (x"c0",x"02",x"9a",x"4a"),
  2866 => (x"c3",x"1e",x"87",x"ec"),
  2867 => (x"fd",x"49",x"d4",x"c2"),
  2868 => (x"c4",x"87",x"da",x"ee"),
  2869 => (x"02",x"98",x"70",x"86"),
  2870 => (x"f5",x"c2",x"87",x"dc"),
  2871 => (x"c2",x"c3",x"1e",x"de"),
  2872 => (x"f1",x"fd",x"49",x"d4"),
  2873 => (x"86",x"c4",x"87",x"dc"),
  2874 => (x"c9",x"02",x"98",x"70"),
  2875 => (x"de",x"f5",x"c2",x"87"),
  2876 => (x"87",x"dd",x"fe",x"49"),
  2877 => (x"48",x"c0",x"87",x"c2"),
  2878 => (x"71",x"1e",x"4f",x"26"),
  2879 => (x"c0",x"02",x"9a",x"4a"),
  2880 => (x"c3",x"1e",x"87",x"ee"),
  2881 => (x"fd",x"49",x"d4",x"c2"),
  2882 => (x"c4",x"87",x"e2",x"ed"),
  2883 => (x"02",x"98",x"70",x"86"),
  2884 => (x"f5",x"c2",x"87",x"de"),
  2885 => (x"d7",x"fe",x"49",x"de"),
  2886 => (x"de",x"f5",x"c2",x"87"),
  2887 => (x"d4",x"c2",x"c3",x"1e"),
  2888 => (x"ec",x"f1",x"fd",x"49"),
  2889 => (x"70",x"86",x"c4",x"87"),
  2890 => (x"87",x"c4",x"02",x"98"),
  2891 => (x"87",x"c2",x"48",x"c1"),
  2892 => (x"4f",x"26",x"48",x"c0"),
  2893 => (x"00",x"00",x"00",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

