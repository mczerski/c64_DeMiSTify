library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"d0c8c387",
    12 => x"86c0c64e",
    13 => x"49d0c8c3",
    14 => x"48f8f4c2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087c3e6",
    19 => x"1e87fc98",
    20 => x"1e731e72",
    21 => x"02114812",
    22 => x"c34b87ca",
    23 => x"739b98df",
    24 => x"87f00288",
    25 => x"4a264b26",
    26 => x"731e4f26",
    27 => x"c11e721e",
    28 => x"87ca048b",
    29 => x"02114812",
    30 => x"028887c4",
    31 => x"4a2687f1",
    32 => x"4f264b26",
    33 => x"731e741e",
    34 => x"c11e721e",
    35 => x"87d0048b",
    36 => x"02114812",
    37 => x"c34c87ca",
    38 => x"749c98df",
    39 => x"87eb0288",
    40 => x"4b264a26",
    41 => x"4f264c26",
    42 => x"8148731e",
    43 => x"c502a973",
    44 => x"05531287",
    45 => x"4f2687f6",
    46 => x"4a66c41e",
    47 => x"51124871",
    48 => x"2687fb05",
    49 => x"4a711e4f",
    50 => x"484966c4",
    51 => x"a6c888c1",
    52 => x"02997158",
    53 => x"481287d4",
    54 => x"7808d4ff",
    55 => x"484966c4",
    56 => x"a6c888c1",
    57 => x"05997158",
    58 => x"4f2687ec",
    59 => x"c44a711e",
    60 => x"c1484966",
    61 => x"58a6c888",
    62 => x"d6029971",
    63 => x"48d4ff87",
    64 => x"6878ffc3",
    65 => x"4966c452",
    66 => x"c888c148",
    67 => x"997158a6",
    68 => x"2687ea05",
    69 => x"1e731e4f",
    70 => x"c34bd4ff",
    71 => x"4a6b7bff",
    72 => x"6b7bffc3",
    73 => x"7232c849",
    74 => x"7bffc3b1",
    75 => x"31c84a6b",
    76 => x"ffc3b271",
    77 => x"c8496b7b",
    78 => x"71b17232",
    79 => x"2687c448",
    80 => x"264c264d",
    81 => x"0e4f264b",
    82 => x"5d5c5b5e",
    83 => x"ff4a710e",
    84 => x"49724cd4",
    85 => x"7199ffc3",
    86 => x"f8f4c27c",
    87 => x"87c805bf",
    88 => x"c94866d0",
    89 => x"58a6d430",
    90 => x"d84966d0",
    91 => x"99ffc329",
    92 => x"66d07c71",
    93 => x"c329d049",
    94 => x"7c7199ff",
    95 => x"c84966d0",
    96 => x"99ffc329",
    97 => x"66d07c71",
    98 => x"99ffc349",
    99 => x"49727c71",
   100 => x"ffc329d0",
   101 => x"6c7c7199",
   102 => x"fff0c94b",
   103 => x"abffc34d",
   104 => x"c387d005",
   105 => x"4b6c7cff",
   106 => x"c6028dc1",
   107 => x"abffc387",
   108 => x"7387f002",
   109 => x"87c7fe48",
   110 => x"ff49c01e",
   111 => x"ffc348d4",
   112 => x"c381c178",
   113 => x"04a9b7c8",
   114 => x"4f2687f1",
   115 => x"e71e731e",
   116 => x"dff8c487",
   117 => x"c01ec04b",
   118 => x"f7c1f0ff",
   119 => x"87e7fd49",
   120 => x"a8c186c4",
   121 => x"87eac005",
   122 => x"c348d4ff",
   123 => x"c0c178ff",
   124 => x"c0c0c0c0",
   125 => x"f0e1c01e",
   126 => x"fd49e9c1",
   127 => x"86c487c9",
   128 => x"ca059870",
   129 => x"48d4ff87",
   130 => x"c178ffc3",
   131 => x"fe87cb48",
   132 => x"8bc187e6",
   133 => x"87fdfe05",
   134 => x"e6fc48c0",
   135 => x"1e731e87",
   136 => x"c348d4ff",
   137 => x"4bd378ff",
   138 => x"ffc01ec0",
   139 => x"49c1c1f0",
   140 => x"c487d4fc",
   141 => x"05987086",
   142 => x"d4ff87ca",
   143 => x"78ffc348",
   144 => x"87cb48c1",
   145 => x"c187f1fd",
   146 => x"dbff058b",
   147 => x"fb48c087",
   148 => x"5e0e87f1",
   149 => x"ff0e5c5b",
   150 => x"dbfd4cd4",
   151 => x"1eeac687",
   152 => x"c1f0e1c0",
   153 => x"defb49c8",
   154 => x"c186c487",
   155 => x"87c802a8",
   156 => x"c087eafe",
   157 => x"87e2c148",
   158 => x"7087dafa",
   159 => x"ffffcf49",
   160 => x"a9eac699",
   161 => x"fe87c802",
   162 => x"48c087d3",
   163 => x"c387cbc1",
   164 => x"f1c07cff",
   165 => x"87f4fc4b",
   166 => x"c0029870",
   167 => x"1ec087eb",
   168 => x"c1f0ffc0",
   169 => x"defa49fa",
   170 => x"7086c487",
   171 => x"87d90598",
   172 => x"6c7cffc3",
   173 => x"7cffc349",
   174 => x"c17c7c7c",
   175 => x"c40299c0",
   176 => x"d548c187",
   177 => x"d148c087",
   178 => x"05abc287",
   179 => x"48c087c4",
   180 => x"8bc187c8",
   181 => x"87fdfe05",
   182 => x"e4f948c0",
   183 => x"1e731e87",
   184 => x"48f8f4c2",
   185 => x"4bc778c1",
   186 => x"c248d0ff",
   187 => x"87c8fb78",
   188 => x"c348d0ff",
   189 => x"c01ec078",
   190 => x"c0c1d0e5",
   191 => x"87c7f949",
   192 => x"a8c186c4",
   193 => x"4b87c105",
   194 => x"c505abc2",
   195 => x"c048c087",
   196 => x"8bc187f9",
   197 => x"87d0ff05",
   198 => x"c287f7fc",
   199 => x"7058fcf4",
   200 => x"87cd0598",
   201 => x"ffc01ec1",
   202 => x"49d0c1f0",
   203 => x"c487d8f8",
   204 => x"48d4ff86",
   205 => x"c478ffc3",
   206 => x"f5c287de",
   207 => x"d0ff58c0",
   208 => x"ff78c248",
   209 => x"ffc348d4",
   210 => x"f748c178",
   211 => x"5e0e87f5",
   212 => x"0e5d5c5b",
   213 => x"ffc34a71",
   214 => x"4cd4ff4d",
   215 => x"d0ff7c75",
   216 => x"78c3c448",
   217 => x"1e727c75",
   218 => x"c1f0ffc0",
   219 => x"d6f749d8",
   220 => x"7086c487",
   221 => x"87c50298",
   222 => x"f0c048c1",
   223 => x"c37c7587",
   224 => x"c0c87cfe",
   225 => x"4966d41e",
   226 => x"c487faf4",
   227 => x"757c7586",
   228 => x"d87c757c",
   229 => x"754be0da",
   230 => x"99496c7c",
   231 => x"c187c505",
   232 => x"87f3058b",
   233 => x"d0ff7c75",
   234 => x"c078c248",
   235 => x"87cff648",
   236 => x"5c5b5e0e",
   237 => x"4b710e5d",
   238 => x"eec54cc0",
   239 => x"ff4adfcd",
   240 => x"ffc348d4",
   241 => x"c3496878",
   242 => x"c005a9fe",
   243 => x"4d7087fd",
   244 => x"cc029b73",
   245 => x"1e66d087",
   246 => x"cff44973",
   247 => x"d686c487",
   248 => x"48d0ff87",
   249 => x"c378d1c4",
   250 => x"66d07dff",
   251 => x"d488c148",
   252 => x"987058a6",
   253 => x"ff87f005",
   254 => x"ffc348d4",
   255 => x"9b737878",
   256 => x"ff87c505",
   257 => x"78d048d0",
   258 => x"c14c4ac1",
   259 => x"eefe058a",
   260 => x"f4487487",
   261 => x"731e87e9",
   262 => x"c04a711e",
   263 => x"48d4ff4b",
   264 => x"ff78ffc3",
   265 => x"c3c448d0",
   266 => x"48d4ff78",
   267 => x"7278ffc3",
   268 => x"f0ffc01e",
   269 => x"f449d1c1",
   270 => x"86c487cd",
   271 => x"d2059870",
   272 => x"1ec0c887",
   273 => x"fd4966cc",
   274 => x"86c487e6",
   275 => x"d0ff4b70",
   276 => x"7378c248",
   277 => x"87ebf348",
   278 => x"5c5b5e0e",
   279 => x"1ec00e5d",
   280 => x"c1f0ffc0",
   281 => x"def349c9",
   282 => x"c21ed287",
   283 => x"fc49c0f5",
   284 => x"86c887fe",
   285 => x"84c14cc0",
   286 => x"04acb7d2",
   287 => x"f5c287f8",
   288 => x"49bf97c0",
   289 => x"c199c0c3",
   290 => x"c005a9c0",
   291 => x"f5c287e7",
   292 => x"49bf97c7",
   293 => x"f5c231d0",
   294 => x"4abf97c8",
   295 => x"b17232c8",
   296 => x"97c9f5c2",
   297 => x"71b14abf",
   298 => x"ffffcf4c",
   299 => x"84c19cff",
   300 => x"e7c134ca",
   301 => x"c9f5c287",
   302 => x"c149bf97",
   303 => x"c299c631",
   304 => x"bf97caf5",
   305 => x"2ab7c74a",
   306 => x"f5c2b172",
   307 => x"4abf97c5",
   308 => x"c29dcf4d",
   309 => x"bf97c6f5",
   310 => x"ca9ac34a",
   311 => x"c7f5c232",
   312 => x"c24bbf97",
   313 => x"c2b27333",
   314 => x"bf97c8f5",
   315 => x"9bc0c34b",
   316 => x"732bb7c6",
   317 => x"c181c2b2",
   318 => x"70307148",
   319 => x"7548c149",
   320 => x"724d7030",
   321 => x"7184c14c",
   322 => x"b7c0c894",
   323 => x"87cc06ad",
   324 => x"2db734c1",
   325 => x"adb7c0c8",
   326 => x"87f4ff01",
   327 => x"def04874",
   328 => x"5b5e0e87",
   329 => x"f80e5d5c",
   330 => x"e6fdc286",
   331 => x"c278c048",
   332 => x"c01edef5",
   333 => x"87defb49",
   334 => x"987086c4",
   335 => x"c087c505",
   336 => x"87cec948",
   337 => x"7ec14dc0",
   338 => x"bfc0f3c0",
   339 => x"d4f6c249",
   340 => x"4bc8714a",
   341 => x"7087d3ec",
   342 => x"87c20598",
   343 => x"f2c07ec0",
   344 => x"c249bffc",
   345 => x"714af0f6",
   346 => x"fdeb4bc8",
   347 => x"05987087",
   348 => x"7ec087c2",
   349 => x"fdc0026e",
   350 => x"e4fcc287",
   351 => x"fdc24dbf",
   352 => x"7ebf9fdc",
   353 => x"ead6c548",
   354 => x"87c705a8",
   355 => x"bfe4fcc2",
   356 => x"6e87ce4d",
   357 => x"d5e9ca48",
   358 => x"87c502a8",
   359 => x"f1c748c0",
   360 => x"def5c287",
   361 => x"f949751e",
   362 => x"86c487ec",
   363 => x"c5059870",
   364 => x"c748c087",
   365 => x"f2c087dc",
   366 => x"c249bffc",
   367 => x"714af0f6",
   368 => x"e5ea4bc8",
   369 => x"05987087",
   370 => x"fdc287c8",
   371 => x"78c148e6",
   372 => x"f3c087da",
   373 => x"c249bfc0",
   374 => x"714ad4f6",
   375 => x"c9ea4bc8",
   376 => x"02987087",
   377 => x"c087c5c0",
   378 => x"87e6c648",
   379 => x"97dcfdc2",
   380 => x"d5c149bf",
   381 => x"cdc005a9",
   382 => x"ddfdc287",
   383 => x"c249bf97",
   384 => x"c002a9ea",
   385 => x"48c087c5",
   386 => x"c287c7c6",
   387 => x"bf97def5",
   388 => x"e9c3487e",
   389 => x"cec002a8",
   390 => x"c3486e87",
   391 => x"c002a8eb",
   392 => x"48c087c5",
   393 => x"c287ebc5",
   394 => x"bf97e9f5",
   395 => x"c0059949",
   396 => x"f5c287cc",
   397 => x"49bf97ea",
   398 => x"c002a9c2",
   399 => x"48c087c5",
   400 => x"c287cfc5",
   401 => x"bf97ebf5",
   402 => x"e2fdc248",
   403 => x"484c7058",
   404 => x"fdc288c1",
   405 => x"f5c258e6",
   406 => x"49bf97ec",
   407 => x"f5c28175",
   408 => x"4abf97ed",
   409 => x"a17232c8",
   410 => x"f3c1c37e",
   411 => x"c2786e48",
   412 => x"bf97eef5",
   413 => x"58a6c848",
   414 => x"bfe6fdc2",
   415 => x"87d4c202",
   416 => x"bffcf2c0",
   417 => x"f0f6c249",
   418 => x"4bc8714a",
   419 => x"7087dbe7",
   420 => x"c5c00298",
   421 => x"c348c087",
   422 => x"fdc287f8",
   423 => x"c34cbfde",
   424 => x"c25cc7c2",
   425 => x"bf97c3f6",
   426 => x"c231c849",
   427 => x"bf97c2f6",
   428 => x"c249a14a",
   429 => x"bf97c4f6",
   430 => x"7232d04a",
   431 => x"f6c249a1",
   432 => x"4abf97c5",
   433 => x"a17232d8",
   434 => x"9166c449",
   435 => x"bff3c1c3",
   436 => x"fbc1c381",
   437 => x"cbf6c259",
   438 => x"c84abf97",
   439 => x"caf6c232",
   440 => x"a24bbf97",
   441 => x"ccf6c24a",
   442 => x"d04bbf97",
   443 => x"4aa27333",
   444 => x"97cdf6c2",
   445 => x"9bcf4bbf",
   446 => x"a27333d8",
   447 => x"ffc1c34a",
   448 => x"fbc1c35a",
   449 => x"8ac24abf",
   450 => x"c1c39274",
   451 => x"a17248ff",
   452 => x"87cac178",
   453 => x"97f0f5c2",
   454 => x"31c849bf",
   455 => x"97eff5c2",
   456 => x"49a14abf",
   457 => x"59eefdc2",
   458 => x"bfeafdc2",
   459 => x"c731c549",
   460 => x"29c981ff",
   461 => x"59c7c2c3",
   462 => x"97f5f5c2",
   463 => x"32c84abf",
   464 => x"97f4f5c2",
   465 => x"4aa24bbf",
   466 => x"6e9266c4",
   467 => x"c3c2c382",
   468 => x"fbc1c35a",
   469 => x"c378c048",
   470 => x"7248f7c1",
   471 => x"c2c378a1",
   472 => x"c1c348c7",
   473 => x"c378bffb",
   474 => x"c348cbc2",
   475 => x"78bfffc1",
   476 => x"bfe6fdc2",
   477 => x"87c9c002",
   478 => x"30c44874",
   479 => x"c9c07e70",
   480 => x"c3c2c387",
   481 => x"30c448bf",
   482 => x"fdc27e70",
   483 => x"786e48ea",
   484 => x"8ef848c1",
   485 => x"4c264d26",
   486 => x"4f264b26",
   487 => x"5c5b5e0e",
   488 => x"4a710e5d",
   489 => x"bfe6fdc2",
   490 => x"7287cb02",
   491 => x"722bc74b",
   492 => x"9cffc14c",
   493 => x"4b7287c9",
   494 => x"4c722bc8",
   495 => x"c39cffc3",
   496 => x"83bff3c1",
   497 => x"bff8f2c0",
   498 => x"87d902ab",
   499 => x"5bfcf2c0",
   500 => x"1edef5c2",
   501 => x"fdf04973",
   502 => x"7086c487",
   503 => x"87c50598",
   504 => x"e6c048c0",
   505 => x"e6fdc287",
   506 => x"87d202bf",
   507 => x"91c44974",
   508 => x"81def5c2",
   509 => x"ffcf4d69",
   510 => x"9dffffff",
   511 => x"497487cb",
   512 => x"f5c291c2",
   513 => x"699f81de",
   514 => x"fe48754d",
   515 => x"5e0e87c6",
   516 => x"0e5d5c5b",
   517 => x"c04d711e",
   518 => x"ca49c11e",
   519 => x"86c487ff",
   520 => x"029c4c70",
   521 => x"c287c0c1",
   522 => x"754aeefd",
   523 => x"87dfe049",
   524 => x"c0029870",
   525 => x"4a7487f1",
   526 => x"4bcb4975",
   527 => x"7087c5e1",
   528 => x"e2c00298",
   529 => x"741ec087",
   530 => x"87c7029c",
   531 => x"c048a6c4",
   532 => x"c487c578",
   533 => x"78c148a6",
   534 => x"c94966c4",
   535 => x"86c487ff",
   536 => x"059c4c70",
   537 => x"7487c0ff",
   538 => x"e7fc2648",
   539 => x"5b5e0e87",
   540 => x"1e0e5d5c",
   541 => x"059b4b71",
   542 => x"48c087c5",
   543 => x"c887e5c1",
   544 => x"7dc04da3",
   545 => x"c70266d4",
   546 => x"9766d487",
   547 => x"87c505bf",
   548 => x"cfc148c0",
   549 => x"4966d487",
   550 => x"7087f3fd",
   551 => x"c1029c4c",
   552 => x"a4dc87c0",
   553 => x"da7d6949",
   554 => x"a3c449a4",
   555 => x"7a699f4a",
   556 => x"bfe6fdc2",
   557 => x"d487d202",
   558 => x"699f49a4",
   559 => x"ffffc049",
   560 => x"d0487199",
   561 => x"c27e7030",
   562 => x"6e7ec087",
   563 => x"806a4849",
   564 => x"7bc07a70",
   565 => x"6a49a3cc",
   566 => x"49a3d079",
   567 => x"48c179c0",
   568 => x"48c087c2",
   569 => x"87ecfa26",
   570 => x"5c5b5e0e",
   571 => x"4c710e5d",
   572 => x"cac1029c",
   573 => x"49a4c887",
   574 => x"c2c10269",
   575 => x"4a66d087",
   576 => x"d482496c",
   577 => x"66d05aa6",
   578 => x"fdc2b94d",
   579 => x"ff4abfe2",
   580 => x"719972ba",
   581 => x"e4c00299",
   582 => x"4ba4c487",
   583 => x"fbf9496b",
   584 => x"c27b7087",
   585 => x"49bfdefd",
   586 => x"7c71816c",
   587 => x"fdc2b975",
   588 => x"ff4abfe2",
   589 => x"719972ba",
   590 => x"dcff0599",
   591 => x"f97c7587",
   592 => x"731e87d2",
   593 => x"9b4b711e",
   594 => x"c887c702",
   595 => x"056949a3",
   596 => x"48c087c5",
   597 => x"c387f7c0",
   598 => x"4abff7c1",
   599 => x"6949a3c4",
   600 => x"c289c249",
   601 => x"91bfdefd",
   602 => x"c24aa271",
   603 => x"49bfe2fd",
   604 => x"a271996b",
   605 => x"fcf2c04a",
   606 => x"1e66c85a",
   607 => x"d5ea4972",
   608 => x"7086c487",
   609 => x"87c40598",
   610 => x"87c248c0",
   611 => x"c7f848c1",
   612 => x"1e731e87",
   613 => x"029b4b71",
   614 => x"a3c887c7",
   615 => x"c5056949",
   616 => x"c048c087",
   617 => x"c1c387f7",
   618 => x"c44abff7",
   619 => x"496949a3",
   620 => x"fdc289c2",
   621 => x"7191bfde",
   622 => x"fdc24aa2",
   623 => x"6b49bfe2",
   624 => x"4aa27199",
   625 => x"5afcf2c0",
   626 => x"721e66c8",
   627 => x"87fee549",
   628 => x"987086c4",
   629 => x"c087c405",
   630 => x"c187c248",
   631 => x"87f8f648",
   632 => x"5c5b5e0e",
   633 => x"711e0e5d",
   634 => x"4c66d44b",
   635 => x"9b732cc9",
   636 => x"87cfc102",
   637 => x"6949a3c8",
   638 => x"87c7c102",
   639 => x"d44da3d0",
   640 => x"fdc27d66",
   641 => x"ff49bfe2",
   642 => x"994a6bb9",
   643 => x"03ac717e",
   644 => x"7bc087cd",
   645 => x"4aa3cc7d",
   646 => x"6a49a3c4",
   647 => x"7287c279",
   648 => x"029c748c",
   649 => x"1e4987dd",
   650 => x"fbfa4973",
   651 => x"d486c487",
   652 => x"ffc74966",
   653 => x"87cb0299",
   654 => x"1edef5c2",
   655 => x"c1fc4973",
   656 => x"2686c487",
   657 => x"1e87cdf5",
   658 => x"4b711e73",
   659 => x"e4c0029b",
   660 => x"cbc2c387",
   661 => x"c24a735b",
   662 => x"defdc28a",
   663 => x"c39249bf",
   664 => x"48bff7c1",
   665 => x"c2c38072",
   666 => x"487158cf",
   667 => x"fdc230c4",
   668 => x"edc058ee",
   669 => x"c7c2c387",
   670 => x"fbc1c348",
   671 => x"c2c378bf",
   672 => x"c1c348cb",
   673 => x"c278bfff",
   674 => x"02bfe6fd",
   675 => x"fdc287c9",
   676 => x"c449bfde",
   677 => x"c387c731",
   678 => x"49bfc3c2",
   679 => x"fdc231c4",
   680 => x"f3f359ee",
   681 => x"5b5e0e87",
   682 => x"4a710e5c",
   683 => x"9a724bc0",
   684 => x"87e1c002",
   685 => x"9f49a2da",
   686 => x"fdc24b69",
   687 => x"cf02bfe6",
   688 => x"49a2d487",
   689 => x"4c49699f",
   690 => x"9cffffc0",
   691 => x"87c234d0",
   692 => x"49744cc0",
   693 => x"fd4973b3",
   694 => x"f9f287ed",
   695 => x"5b5e0e87",
   696 => x"f40e5d5c",
   697 => x"c04a7186",
   698 => x"029a727e",
   699 => x"f5c287d8",
   700 => x"78c048da",
   701 => x"48d2f5c2",
   702 => x"bfcbc2c3",
   703 => x"d6f5c278",
   704 => x"c7c2c348",
   705 => x"fdc278bf",
   706 => x"50c048fb",
   707 => x"bfeafdc2",
   708 => x"daf5c249",
   709 => x"aa714abf",
   710 => x"87c9c403",
   711 => x"99cf4972",
   712 => x"87e9c005",
   713 => x"48f8f2c0",
   714 => x"bfd2f5c2",
   715 => x"def5c278",
   716 => x"d2f5c21e",
   717 => x"f5c249bf",
   718 => x"a1c148d2",
   719 => x"d5e37178",
   720 => x"c086c487",
   721 => x"c248f4f2",
   722 => x"cc78def5",
   723 => x"f4f2c087",
   724 => x"e0c048bf",
   725 => x"f8f2c080",
   726 => x"daf5c258",
   727 => x"80c148bf",
   728 => x"58def5c2",
   729 => x"000cb427",
   730 => x"bf97bf00",
   731 => x"c2029d4d",
   732 => x"e5c387e3",
   733 => x"dcc202ad",
   734 => x"f4f2c087",
   735 => x"a3cb4bbf",
   736 => x"cf4c1149",
   737 => x"d2c105ac",
   738 => x"df497587",
   739 => x"cd89c199",
   740 => x"eefdc291",
   741 => x"4aa3c181",
   742 => x"a3c35112",
   743 => x"c551124a",
   744 => x"51124aa3",
   745 => x"124aa3c7",
   746 => x"4aa3c951",
   747 => x"a3ce5112",
   748 => x"d051124a",
   749 => x"51124aa3",
   750 => x"124aa3d2",
   751 => x"4aa3d451",
   752 => x"a3d65112",
   753 => x"d851124a",
   754 => x"51124aa3",
   755 => x"124aa3dc",
   756 => x"4aa3de51",
   757 => x"7ec15112",
   758 => x"7487fac0",
   759 => x"0599c849",
   760 => x"7487ebc0",
   761 => x"0599d049",
   762 => x"66dc87d1",
   763 => x"87cbc002",
   764 => x"66dc4973",
   765 => x"0298700f",
   766 => x"6e87d3c0",
   767 => x"87c6c005",
   768 => x"48eefdc2",
   769 => x"f2c050c0",
   770 => x"c248bff4",
   771 => x"fdc287e1",
   772 => x"50c048fb",
   773 => x"eafdc27e",
   774 => x"f5c249bf",
   775 => x"714abfda",
   776 => x"f7fb04aa",
   777 => x"cbc2c387",
   778 => x"c8c005bf",
   779 => x"e6fdc287",
   780 => x"f8c102bf",
   781 => x"d6f5c287",
   782 => x"dfed49bf",
   783 => x"c2497087",
   784 => x"c459daf5",
   785 => x"f5c248a6",
   786 => x"c278bfd6",
   787 => x"02bfe6fd",
   788 => x"c487d8c0",
   789 => x"ffcf4966",
   790 => x"99f8ffff",
   791 => x"c5c002a9",
   792 => x"c04cc087",
   793 => x"4cc187e1",
   794 => x"c487dcc0",
   795 => x"ffcf4966",
   796 => x"02a999f8",
   797 => x"c887c8c0",
   798 => x"78c048a6",
   799 => x"c887c5c0",
   800 => x"78c148a6",
   801 => x"744c66c8",
   802 => x"e0c0059c",
   803 => x"4966c487",
   804 => x"fdc289c2",
   805 => x"914abfde",
   806 => x"bff7c1c3",
   807 => x"d2f5c24a",
   808 => x"78a17248",
   809 => x"48daf5c2",
   810 => x"dff978c0",
   811 => x"f448c087",
   812 => x"87e0eb8e",
   813 => x"00000000",
   814 => x"ffffffff",
   815 => x"00000cc4",
   816 => x"00000ccd",
   817 => x"33544146",
   818 => x"20202032",
   819 => x"54414600",
   820 => x"20203631",
   821 => x"ff1e0020",
   822 => x"ffc348d4",
   823 => x"26486878",
   824 => x"d4ff1e4f",
   825 => x"78ffc348",
   826 => x"c848d0ff",
   827 => x"d4ff78e1",
   828 => x"c378d448",
   829 => x"ff48cfc2",
   830 => x"2650bfd4",
   831 => x"d0ff1e4f",
   832 => x"78e0c048",
   833 => x"ff1e4f26",
   834 => x"497087cc",
   835 => x"87c60299",
   836 => x"05a9fbc0",
   837 => x"487187f1",
   838 => x"5e0e4f26",
   839 => x"710e5c5b",
   840 => x"fe4cc04b",
   841 => x"497087f0",
   842 => x"f9c00299",
   843 => x"a9ecc087",
   844 => x"87f2c002",
   845 => x"02a9fbc0",
   846 => x"cc87ebc0",
   847 => x"03acb766",
   848 => x"66d087c7",
   849 => x"7187c202",
   850 => x"02997153",
   851 => x"84c187c2",
   852 => x"7087c3fe",
   853 => x"cd029949",
   854 => x"a9ecc087",
   855 => x"c087c702",
   856 => x"ff05a9fb",
   857 => x"66d087d5",
   858 => x"c087c302",
   859 => x"ecc07b97",
   860 => x"87c405a9",
   861 => x"87c54a74",
   862 => x"0ac04a74",
   863 => x"c248728a",
   864 => x"264d2687",
   865 => x"264b264c",
   866 => x"c9fd1e4f",
   867 => x"c0497087",
   868 => x"04a9b7f0",
   869 => x"f9c087ca",
   870 => x"c301a9b7",
   871 => x"89f0c087",
   872 => x"a9b7c1c1",
   873 => x"c187ca04",
   874 => x"01a9b7da",
   875 => x"f7c087c3",
   876 => x"b7e1c189",
   877 => x"87ca04a9",
   878 => x"a9b7fac1",
   879 => x"c087c301",
   880 => x"487189fd",
   881 => x"5e0e4f26",
   882 => x"710e5c5b",
   883 => x"4cd4ff4a",
   884 => x"eac04972",
   885 => x"9b4b7087",
   886 => x"c187c202",
   887 => x"48d0ff8b",
   888 => x"c178c5c8",
   889 => x"49737cd5",
   890 => x"e7c131c6",
   891 => x"4abf97e5",
   892 => x"70b07148",
   893 => x"48d0ff7c",
   894 => x"487378c4",
   895 => x"0e87c4fe",
   896 => x"5d5c5b5e",
   897 => x"7186f80e",
   898 => x"c07ec04b",
   899 => x"bf97e6fb",
   900 => x"05a9df49",
   901 => x"c887eec0",
   902 => x"699749a3",
   903 => x"a9c3c149",
   904 => x"c987dd05",
   905 => x"699749a3",
   906 => x"a9c6c149",
   907 => x"ca87d105",
   908 => x"699749a3",
   909 => x"a9c7c149",
   910 => x"c187c505",
   911 => x"87e1c248",
   912 => x"dcc248c0",
   913 => x"87d9fa87",
   914 => x"fbc04cc0",
   915 => x"49bf97e6",
   916 => x"cf04a9c0",
   917 => x"87eefa87",
   918 => x"fbc084c1",
   919 => x"49bf97e6",
   920 => x"87f106ac",
   921 => x"97e6fbc0",
   922 => x"87cf02bf",
   923 => x"7087e7f9",
   924 => x"c6029949",
   925 => x"a9ecc087",
   926 => x"c087f105",
   927 => x"87d6f94c",
   928 => x"d1f94d70",
   929 => x"58a6c887",
   930 => x"7087cbf9",
   931 => x"c884c14a",
   932 => x"699749a3",
   933 => x"c702ad49",
   934 => x"adffc087",
   935 => x"87e7c005",
   936 => x"9749a3c9",
   937 => x"66c44969",
   938 => x"87c702a9",
   939 => x"a8ffc048",
   940 => x"ca87d405",
   941 => x"699749a3",
   942 => x"c602aa49",
   943 => x"aaffc087",
   944 => x"c187c405",
   945 => x"c087d07e",
   946 => x"c602adec",
   947 => x"adfbc087",
   948 => x"c087c405",
   949 => x"6e7ec14c",
   950 => x"87e1fe02",
   951 => x"7487def8",
   952 => x"fa8ef848",
   953 => x"0e0087db",
   954 => x"5d5c5b5e",
   955 => x"4d711e0e",
   956 => x"754bd4ff",
   957 => x"d4c2c31e",
   958 => x"87f1e549",
   959 => x"987086c4",
   960 => x"87d8c302",
   961 => x"bfdcc2c3",
   962 => x"fa49754c",
   963 => x"d0ff87f8",
   964 => x"78c5c848",
   965 => x"c07bd6c1",
   966 => x"49a2754a",
   967 => x"82c17b11",
   968 => x"04aab7cb",
   969 => x"4acc87f3",
   970 => x"c17bffc3",
   971 => x"b7e0c082",
   972 => x"87f404aa",
   973 => x"c448d0ff",
   974 => x"7bffc378",
   975 => x"c178c5c8",
   976 => x"7bc17bd3",
   977 => x"9c7478c4",
   978 => x"87ffc102",
   979 => x"7edef5c2",
   980 => x"8c4dc0c8",
   981 => x"03acb7c0",
   982 => x"c0c887c6",
   983 => x"4cc04da4",
   984 => x"05adc0c8",
   985 => x"c2c387dc",
   986 => x"49bf97cf",
   987 => x"d10299d0",
   988 => x"c31ec087",
   989 => x"e749d4c2",
   990 => x"86c487c8",
   991 => x"c04a4970",
   992 => x"f5c287ee",
   993 => x"c2c31ede",
   994 => x"f5e649d4",
   995 => x"7086c487",
   996 => x"d0ff4a49",
   997 => x"78c5c848",
   998 => x"6e7bd4c1",
   999 => x"6e7bbf97",
  1000 => x"7080c148",
  1001 => x"058dc17e",
  1002 => x"ff87f0ff",
  1003 => x"78c448d0",
  1004 => x"c5059a72",
  1005 => x"c048c087",
  1006 => x"1ec187e4",
  1007 => x"49d4c2c3",
  1008 => x"c487e5e4",
  1009 => x"059c7486",
  1010 => x"ff87c1fe",
  1011 => x"c5c848d0",
  1012 => x"7bd3c178",
  1013 => x"78c47bc0",
  1014 => x"87c248c1",
  1015 => x"262648c0",
  1016 => x"264c264d",
  1017 => x"0e4f264b",
  1018 => x"5d5c5b5e",
  1019 => x"4b711e0e",
  1020 => x"ab4d4cc0",
  1021 => x"87e8c004",
  1022 => x"1efff7c0",
  1023 => x"c4029d75",
  1024 => x"c24ac087",
  1025 => x"724ac187",
  1026 => x"87d1eb49",
  1027 => x"7e7086c4",
  1028 => x"056e84c1",
  1029 => x"4c7387c2",
  1030 => x"ac7385c1",
  1031 => x"87d8ff06",
  1032 => x"fe26486e",
  1033 => x"5e0e87f9",
  1034 => x"710e5c5b",
  1035 => x"0266cc4b",
  1036 => x"4c87e8c0",
  1037 => x"028cf0c0",
  1038 => x"7487e8c0",
  1039 => x"028ac14a",
  1040 => x"8a87e0c0",
  1041 => x"8a87dc02",
  1042 => x"c087d802",
  1043 => x"c0028ae0",
  1044 => x"8ac187e5",
  1045 => x"87e7c002",
  1046 => x"7387eac0",
  1047 => x"87c7fa49",
  1048 => x"7487e2c0",
  1049 => x"c149c01e",
  1050 => x"7487d7ed",
  1051 => x"c149731e",
  1052 => x"c887cfed",
  1053 => x"7387ce86",
  1054 => x"c5f1c149",
  1055 => x"7387c687",
  1056 => x"f5f1c149",
  1057 => x"87d9fd87",
  1058 => x"5c5b5e0e",
  1059 => x"711e0e5d",
  1060 => x"91de494c",
  1061 => x"4dfcc2c3",
  1062 => x"6d978571",
  1063 => x"87dcc102",
  1064 => x"bfe8c2c3",
  1065 => x"7282744a",
  1066 => x"87fbfc49",
  1067 => x"026e7e70",
  1068 => x"c387f2c0",
  1069 => x"6e4bf0c2",
  1070 => x"fe49cb4a",
  1071 => x"7487e9ff",
  1072 => x"c193cb4b",
  1073 => x"c483d8e8",
  1074 => x"c0c4c183",
  1075 => x"c149747b",
  1076 => x"7587fad6",
  1077 => x"e6e7c17b",
  1078 => x"1e49bf97",
  1079 => x"49f0c2c3",
  1080 => x"c487c3fd",
  1081 => x"c1497486",
  1082 => x"c087e2d6",
  1083 => x"c1d8c149",
  1084 => x"d0c2c387",
  1085 => x"c178c048",
  1086 => x"87f0df49",
  1087 => x"87dffb26",
  1088 => x"64616f4c",
  1089 => x"2e676e69",
  1090 => x"0e002e2e",
  1091 => x"0e5c5b5e",
  1092 => x"c34a4b71",
  1093 => x"82bfe8c2",
  1094 => x"cafb4972",
  1095 => x"9c4c7087",
  1096 => x"4987c402",
  1097 => x"c387fee5",
  1098 => x"c048e8c2",
  1099 => x"de49c178",
  1100 => x"ecfa87fa",
  1101 => x"5b5e0e87",
  1102 => x"f40e5d5c",
  1103 => x"def5c286",
  1104 => x"c44cc04d",
  1105 => x"78c048a6",
  1106 => x"bfe8c2c3",
  1107 => x"06a9c049",
  1108 => x"c287c1c1",
  1109 => x"9848def5",
  1110 => x"87f8c002",
  1111 => x"1efff7c0",
  1112 => x"c70266c8",
  1113 => x"48a6c487",
  1114 => x"87c578c0",
  1115 => x"c148a6c4",
  1116 => x"4966c478",
  1117 => x"c487e6e5",
  1118 => x"c14d7086",
  1119 => x"4866c484",
  1120 => x"a6c880c1",
  1121 => x"e8c2c358",
  1122 => x"03ac49bf",
  1123 => x"9d7587c6",
  1124 => x"87c8ff05",
  1125 => x"9d754cc0",
  1126 => x"87e0c302",
  1127 => x"1efff7c0",
  1128 => x"c70266c8",
  1129 => x"48a6cc87",
  1130 => x"87c578c0",
  1131 => x"c148a6cc",
  1132 => x"4966cc78",
  1133 => x"c487e6e4",
  1134 => x"6e7e7086",
  1135 => x"87e9c202",
  1136 => x"81cb496e",
  1137 => x"d0496997",
  1138 => x"d6c10299",
  1139 => x"cbc4c187",
  1140 => x"cb49744a",
  1141 => x"d8e8c191",
  1142 => x"c8797281",
  1143 => x"51ffc381",
  1144 => x"91de4974",
  1145 => x"4dfcc2c3",
  1146 => x"c1c28571",
  1147 => x"a5c17d97",
  1148 => x"51e0c049",
  1149 => x"97eefdc2",
  1150 => x"87d202bf",
  1151 => x"a5c284c1",
  1152 => x"eefdc24b",
  1153 => x"fe49db4a",
  1154 => x"c187ddfa",
  1155 => x"a5cd87db",
  1156 => x"c151c049",
  1157 => x"4ba5c284",
  1158 => x"49cb4a6e",
  1159 => x"87c8fafe",
  1160 => x"c187c6c1",
  1161 => x"744ac8c2",
  1162 => x"c191cb49",
  1163 => x"7281d8e8",
  1164 => x"eefdc279",
  1165 => x"d802bf97",
  1166 => x"de497487",
  1167 => x"c384c191",
  1168 => x"714bfcc2",
  1169 => x"eefdc283",
  1170 => x"fe49dd4a",
  1171 => x"d887d9f9",
  1172 => x"de4b7487",
  1173 => x"fcc2c393",
  1174 => x"49a3cb83",
  1175 => x"84c151c0",
  1176 => x"cb4a6e73",
  1177 => x"fff8fe49",
  1178 => x"4866c487",
  1179 => x"a6c880c1",
  1180 => x"03acc758",
  1181 => x"6e87c5c0",
  1182 => x"87e0fc05",
  1183 => x"8ef44874",
  1184 => x"1e87dcf5",
  1185 => x"4b711e73",
  1186 => x"c191cb49",
  1187 => x"c881d8e8",
  1188 => x"e7c14aa1",
  1189 => x"501248e5",
  1190 => x"c04aa1c9",
  1191 => x"1248e6fb",
  1192 => x"c181ca50",
  1193 => x"1148e6e7",
  1194 => x"e6e7c150",
  1195 => x"1e49bf97",
  1196 => x"f1f549c0",
  1197 => x"d0c2c387",
  1198 => x"c178de48",
  1199 => x"87ecd849",
  1200 => x"87dff426",
  1201 => x"494a711e",
  1202 => x"e8c191cb",
  1203 => x"81c881d8",
  1204 => x"c2c34811",
  1205 => x"c2c358d4",
  1206 => x"78c048e8",
  1207 => x"cbd849c1",
  1208 => x"1e4f2687",
  1209 => x"d0c149c0",
  1210 => x"4f2687c8",
  1211 => x"0299711e",
  1212 => x"e9c187d2",
  1213 => x"50c048ed",
  1214 => x"cbc180f7",
  1215 => x"e8c140c4",
  1216 => x"87ce78c6",
  1217 => x"48e9e9c1",
  1218 => x"78e7e7c1",
  1219 => x"cbc180fc",
  1220 => x"4f2678e3",
  1221 => x"5c5b5e0e",
  1222 => x"4a4c710e",
  1223 => x"e8c192cb",
  1224 => x"a2c882d8",
  1225 => x"4ba2c949",
  1226 => x"1e4b6b97",
  1227 => x"1e496997",
  1228 => x"491282ca",
  1229 => x"87c1f9c0",
  1230 => x"efd649c0",
  1231 => x"c1497487",
  1232 => x"f887cacd",
  1233 => x"87d9f28e",
  1234 => x"711e731e",
  1235 => x"c3ff494b",
  1236 => x"fe497387",
  1237 => x"caf287fe",
  1238 => x"1e731e87",
  1239 => x"a3c64b71",
  1240 => x"87dc024a",
  1241 => x"c0028ac1",
  1242 => x"028a87e4",
  1243 => x"8a87e8c1",
  1244 => x"87cac102",
  1245 => x"efc0028a",
  1246 => x"d9028a87",
  1247 => x"87e9c187",
  1248 => x"48d0c2c3",
  1249 => x"49c178df",
  1250 => x"c187e1d5",
  1251 => x"49c787e6",
  1252 => x"c187f1fc",
  1253 => x"c2c387de",
  1254 => x"c102bfe8",
  1255 => x"c14887cb",
  1256 => x"ecc2c388",
  1257 => x"87c1c158",
  1258 => x"bfecc2c3",
  1259 => x"87f9c002",
  1260 => x"bfe8c2c3",
  1261 => x"c380c148",
  1262 => x"c058ecc2",
  1263 => x"c2c387eb",
  1264 => x"c649bfe8",
  1265 => x"ecc2c389",
  1266 => x"a9b7c059",
  1267 => x"c387da03",
  1268 => x"c048e8c2",
  1269 => x"c387d278",
  1270 => x"02bfecc2",
  1271 => x"c2c387cb",
  1272 => x"c648bfe8",
  1273 => x"ecc2c380",
  1274 => x"d349c058",
  1275 => x"497387fe",
  1276 => x"87d9cac1",
  1277 => x"0e87ecef",
  1278 => x"0e5c5b5e",
  1279 => x"66cc4c71",
  1280 => x"cb4b741e",
  1281 => x"d8e8c193",
  1282 => x"4aa3c483",
  1283 => x"f2fe496a",
  1284 => x"cac187e6",
  1285 => x"a3c87bc3",
  1286 => x"5166d449",
  1287 => x"d849a3c9",
  1288 => x"a3ca5166",
  1289 => x"5166dc49",
  1290 => x"87f5ee26",
  1291 => x"5c5b5e0e",
  1292 => x"d0ff0e5d",
  1293 => x"59a6d886",
  1294 => x"c048a6c8",
  1295 => x"c180fc78",
  1296 => x"c87866c4",
  1297 => x"c478c180",
  1298 => x"c378c180",
  1299 => x"c148ecc2",
  1300 => x"d0c2c378",
  1301 => x"486e7ebf",
  1302 => x"cb05a8de",
  1303 => x"87d5f387",
  1304 => x"a6cc4970",
  1305 => x"87ecd059",
  1306 => x"a8df486e",
  1307 => x"87eec105",
  1308 => x"4966c0c1",
  1309 => x"7e6981c4",
  1310 => x"48c9e3c1",
  1311 => x"a1d0496e",
  1312 => x"7141204a",
  1313 => x"87f905aa",
  1314 => x"4ac3cac1",
  1315 => x"0a66c0c1",
  1316 => x"c0c10a7a",
  1317 => x"81c94966",
  1318 => x"c0c151df",
  1319 => x"81ca4966",
  1320 => x"c151d3c1",
  1321 => x"cb4966c0",
  1322 => x"4ba1c481",
  1323 => x"6b48a6c4",
  1324 => x"721e7178",
  1325 => x"d9e3c11e",
  1326 => x"4966cc48",
  1327 => x"204aa1d0",
  1328 => x"05aa7141",
  1329 => x"4a2687f9",
  1330 => x"79724926",
  1331 => x"df4aa1c9",
  1332 => x"c181ca52",
  1333 => x"a6c851d4",
  1334 => x"ce78c248",
  1335 => x"c0e087f6",
  1336 => x"87e2e087",
  1337 => x"87eedfff",
  1338 => x"fbc04c70",
  1339 => x"d2c102ac",
  1340 => x"0566d487",
  1341 => x"c087c3c1",
  1342 => x"1ec11e1e",
  1343 => x"1ecbeac1",
  1344 => x"f2fb49c0",
  1345 => x"66d0c187",
  1346 => x"6a82c44a",
  1347 => x"7481c749",
  1348 => x"d81ec151",
  1349 => x"c8496a1e",
  1350 => x"fddfff81",
  1351 => x"c186d887",
  1352 => x"c04866c4",
  1353 => x"87c701a8",
  1354 => x"c148a6c8",
  1355 => x"c187cf78",
  1356 => x"c14866c4",
  1357 => x"58a6c888",
  1358 => x"dfff87c4",
  1359 => x"a6cc87c8",
  1360 => x"7478c248",
  1361 => x"c7cd029c",
  1362 => x"4866c887",
  1363 => x"a866c8c1",
  1364 => x"87fccc03",
  1365 => x"c048a6d8",
  1366 => x"c080c478",
  1367 => x"f5ddff78",
  1368 => x"c14c7087",
  1369 => x"c205acd0",
  1370 => x"66dc87db",
  1371 => x"87d9e07e",
  1372 => x"e0c04970",
  1373 => x"ddff59a6",
  1374 => x"4c7087dc",
  1375 => x"05acecc0",
  1376 => x"c887edc1",
  1377 => x"91cb4966",
  1378 => x"8166c0c1",
  1379 => x"6a4aa1c4",
  1380 => x"4aa1c84d",
  1381 => x"c15266dc",
  1382 => x"ff79c4cb",
  1383 => x"7087f7dc",
  1384 => x"d9029c4c",
  1385 => x"acfbc087",
  1386 => x"7487d302",
  1387 => x"e5dcff55",
  1388 => x"9c4c7087",
  1389 => x"c087c702",
  1390 => x"ff05acfb",
  1391 => x"e0c087ed",
  1392 => x"55c1c255",
  1393 => x"d47d97c0",
  1394 => x"a96e4966",
  1395 => x"c887db05",
  1396 => x"66c44866",
  1397 => x"87ca04a8",
  1398 => x"c14866c8",
  1399 => x"58a6cc80",
  1400 => x"66c487c8",
  1401 => x"c888c148",
  1402 => x"dbff58a6",
  1403 => x"4c7087e8",
  1404 => x"05acd0c1",
  1405 => x"66d087c8",
  1406 => x"d480c148",
  1407 => x"d0c158a6",
  1408 => x"e5fd02ac",
  1409 => x"a6e0c087",
  1410 => x"7866d448",
  1411 => x"c04866dc",
  1412 => x"05a866e0",
  1413 => x"c087cbc9",
  1414 => x"c048a6e4",
  1415 => x"48747e78",
  1416 => x"c088fbc0",
  1417 => x"7058a6ec",
  1418 => x"d0c80298",
  1419 => x"88cb4887",
  1420 => x"58a6ecc0",
  1421 => x"c1029870",
  1422 => x"c94887d3",
  1423 => x"a6ecc088",
  1424 => x"02987058",
  1425 => x"4887ddc3",
  1426 => x"ecc088c4",
  1427 => x"987058a6",
  1428 => x"4887d002",
  1429 => x"ecc088c1",
  1430 => x"987058a6",
  1431 => x"87c4c302",
  1432 => x"d887d4c7",
  1433 => x"f0c048a6",
  1434 => x"e9d9ff78",
  1435 => x"c04c7087",
  1436 => x"c002acec",
  1437 => x"a6dc87c3",
  1438 => x"acecc05c",
  1439 => x"87cdc002",
  1440 => x"87d2d9ff",
  1441 => x"ecc04c70",
  1442 => x"f3ff05ac",
  1443 => x"acecc087",
  1444 => x"87c4c002",
  1445 => x"87fed8ff",
  1446 => x"d41e66d8",
  1447 => x"d41e4966",
  1448 => x"c11e4966",
  1449 => x"d81ecbea",
  1450 => x"caf54966",
  1451 => x"ca1ec087",
  1452 => x"66e0c01e",
  1453 => x"c191cb49",
  1454 => x"d88166d8",
  1455 => x"a1c448a6",
  1456 => x"bf66d878",
  1457 => x"d1d9ff49",
  1458 => x"c086d887",
  1459 => x"c106a8b7",
  1460 => x"1ec187c5",
  1461 => x"66c81ede",
  1462 => x"d8ff49bf",
  1463 => x"86c887fc",
  1464 => x"c0484970",
  1465 => x"a6dc8808",
  1466 => x"a8b7c058",
  1467 => x"87e7c006",
  1468 => x"dd4866d8",
  1469 => x"de03a8b7",
  1470 => x"49bf6e87",
  1471 => x"c08166d8",
  1472 => x"66d851e0",
  1473 => x"6e81c149",
  1474 => x"c1c281bf",
  1475 => x"4966d851",
  1476 => x"bf6e81c2",
  1477 => x"cc51c081",
  1478 => x"80c14866",
  1479 => x"c158a6d0",
  1480 => x"87d9c47e",
  1481 => x"87e1d9ff",
  1482 => x"ff58a6dc",
  1483 => x"c087dad9",
  1484 => x"c058a6ec",
  1485 => x"c005a8ec",
  1486 => x"e8c087ca",
  1487 => x"66d848a6",
  1488 => x"87c4c078",
  1489 => x"87ced6ff",
  1490 => x"cb4966c8",
  1491 => x"66c0c191",
  1492 => x"70807148",
  1493 => x"c8496e7e",
  1494 => x"ca4a6e81",
  1495 => x"5266d882",
  1496 => x"4a66e8c0",
  1497 => x"66d882c1",
  1498 => x"7248c18a",
  1499 => x"c14a7030",
  1500 => x"7997728a",
  1501 => x"1e496997",
  1502 => x"c04966dc",
  1503 => x"c487fce6",
  1504 => x"a6f0c086",
  1505 => x"c4496e58",
  1506 => x"c04d6981",
  1507 => x"dc4866e0",
  1508 => x"c002a866",
  1509 => x"a6d887c8",
  1510 => x"c078c048",
  1511 => x"a6d887c5",
  1512 => x"d878c148",
  1513 => x"e0c01e66",
  1514 => x"ff49751e",
  1515 => x"c887ebd5",
  1516 => x"c04c7086",
  1517 => x"c106acb7",
  1518 => x"857487d4",
  1519 => x"7449e0c0",
  1520 => x"c14b7589",
  1521 => x"714ae9e3",
  1522 => x"87dce3fe",
  1523 => x"e4c085c2",
  1524 => x"80c14866",
  1525 => x"58a6e8c0",
  1526 => x"4966ecc0",
  1527 => x"a97081c1",
  1528 => x"87c8c002",
  1529 => x"c048a6d8",
  1530 => x"87c5c078",
  1531 => x"c148a6d8",
  1532 => x"1e66d878",
  1533 => x"c049a4c2",
  1534 => x"887148e0",
  1535 => x"751e4970",
  1536 => x"d5d4ff49",
  1537 => x"c086c887",
  1538 => x"ff01a8b7",
  1539 => x"e4c087c0",
  1540 => x"d1c00266",
  1541 => x"c9496e87",
  1542 => x"66e4c081",
  1543 => x"c1486e51",
  1544 => x"c078d4cc",
  1545 => x"496e87cc",
  1546 => x"51c281c9",
  1547 => x"cdc1486e",
  1548 => x"7ec178c8",
  1549 => x"ff87c6c0",
  1550 => x"7087cbd3",
  1551 => x"c0026e4c",
  1552 => x"66c887f5",
  1553 => x"a866c448",
  1554 => x"87cbc004",
  1555 => x"c14866c8",
  1556 => x"58a6cc80",
  1557 => x"c487e0c0",
  1558 => x"88c14866",
  1559 => x"c058a6c8",
  1560 => x"c6c187d5",
  1561 => x"c8c005ac",
  1562 => x"4866cc87",
  1563 => x"a6d080c1",
  1564 => x"d1d2ff58",
  1565 => x"d04c7087",
  1566 => x"80c14866",
  1567 => x"7458a6d4",
  1568 => x"cbc0029c",
  1569 => x"4866c887",
  1570 => x"a866c8c1",
  1571 => x"87c4f304",
  1572 => x"87e9d1ff",
  1573 => x"c74866c8",
  1574 => x"e5c003a8",
  1575 => x"ecc2c387",
  1576 => x"c878c048",
  1577 => x"91cb4966",
  1578 => x"8166c0c1",
  1579 => x"6a4aa1c4",
  1580 => x"7952c04a",
  1581 => x"c14866c8",
  1582 => x"58a6cc80",
  1583 => x"ff04a8c7",
  1584 => x"d0ff87db",
  1585 => x"d6dcff8e",
  1586 => x"616f4c87",
  1587 => x"65532064",
  1588 => x"6e697474",
  1589 => x"81207367",
  1590 => x"76615300",
  1591 => x"65532065",
  1592 => x"6e697474",
  1593 => x"81207367",
  1594 => x"00203a00",
  1595 => x"711e731e",
  1596 => x"c6029b4b",
  1597 => x"e8c2c387",
  1598 => x"c778c048",
  1599 => x"e8c2c31e",
  1600 => x"c11e49bf",
  1601 => x"c31ed8e8",
  1602 => x"49bfd0c2",
  1603 => x"cc87ddec",
  1604 => x"d0c2c386",
  1605 => x"d3e749bf",
  1606 => x"029b7387",
  1607 => x"e8c187c8",
  1608 => x"f6c049d8",
  1609 => x"daff87f9",
  1610 => x"c11e87f9",
  1611 => x"c149c6e5",
  1612 => x"c187cfce",
  1613 => x"c048e5e7",
  1614 => x"fbe9c150",
  1615 => x"d6ff49bf",
  1616 => x"48c087e5",
  1617 => x"4f434f26",
  1618 => x"20204552",
  1619 => x"46432020",
  1620 => x"ce1e0047",
  1621 => x"49c187c8",
  1622 => x"fe87d1fe",
  1623 => x"7087fee5",
  1624 => x"87cd0298",
  1625 => x"87f9eefe",
  1626 => x"c4029870",
  1627 => x"c24ac187",
  1628 => x"724ac087",
  1629 => x"87ce059a",
  1630 => x"e6c11ec0",
  1631 => x"c1c149e6",
  1632 => x"86c487fa",
  1633 => x"cbc187fe",
  1634 => x"1ec087e2",
  1635 => x"49f1e6c1",
  1636 => x"87e8c1c1",
  1637 => x"d1fe1ec0",
  1638 => x"c1497087",
  1639 => x"c487ddc1",
  1640 => x"8ef887c7",
  1641 => x"44534f26",
  1642 => x"69616620",
  1643 => x"2e64656c",
  1644 => x"6f6f4200",
  1645 => x"676e6974",
  1646 => x"002e2e2e",
  1647 => x"d449c01e",
  1648 => x"f8c087e2",
  1649 => x"c4c187f9",
  1650 => x"87f187e8",
  1651 => x"c31e4f26",
  1652 => x"c048e8c2",
  1653 => x"d0c2c378",
  1654 => x"fd78c048",
  1655 => x"dbff87f4",
  1656 => x"2648c087",
  1657 => x"2000004f",
  1658 => x"20202020",
  1659 => x"20202020",
  1660 => x"20202020",
  1661 => x"74697845",
  1662 => x"20202020",
  1663 => x"20202020",
  1664 => x"20202020",
  1665 => x"20800081",
  1666 => x"20202020",
  1667 => x"20202020",
  1668 => x"42202020",
  1669 => x"006b6361",
  1670 => x"000012c4",
  1671 => x"000030bc",
  1672 => x"c4000000",
  1673 => x"da000012",
  1674 => x"00000030",
  1675 => x"12c40000",
  1676 => x"30f80000",
  1677 => x"00000000",
  1678 => x"0012c400",
  1679 => x"00311600",
  1680 => x"00000000",
  1681 => x"000012c4",
  1682 => x"00003134",
  1683 => x"c4000000",
  1684 => x"52000012",
  1685 => x"00000031",
  1686 => x"12c40000",
  1687 => x"31700000",
  1688 => x"00000000",
  1689 => x"0012c400",
  1690 => x"00000000",
  1691 => x"00000000",
  1692 => x"00001359",
  1693 => x"00000000",
  1694 => x"7f000000",
  1695 => x"4300001a",
  1696 => x"20203436",
  1697 => x"52202020",
  1698 => x"4c004d4f",
  1699 => x"2064616f",
  1700 => x"1e002e2a",
  1701 => x"c048f0fe",
  1702 => x"7909cd78",
  1703 => x"1e4f2609",
  1704 => x"bff0fe1e",
  1705 => x"2626487e",
  1706 => x"f0fe1e4f",
  1707 => x"2678c148",
  1708 => x"f0fe1e4f",
  1709 => x"2678c048",
  1710 => x"4a711e4f",
  1711 => x"c17a97c0",
  1712 => x"51c049a2",
  1713 => x"c049a2ca",
  1714 => x"49a2cb51",
  1715 => x"4f2651c0",
  1716 => x"5c5b5e0e",
  1717 => x"7186f00e",
  1718 => x"49a4ca4c",
  1719 => x"cb7e6997",
  1720 => x"6b974ba4",
  1721 => x"58a6c848",
  1722 => x"a6cc80c1",
  1723 => x"d098c758",
  1724 => x"486e58a6",
  1725 => x"05a866cc",
  1726 => x"699787db",
  1727 => x"486b977e",
  1728 => x"c158a6c8",
  1729 => x"58a6cc80",
  1730 => x"a6d098c7",
  1731 => x"cc486e58",
  1732 => x"e502a866",
  1733 => x"87d9fe87",
  1734 => x"974aa4cc",
  1735 => x"a172496b",
  1736 => x"5166dc49",
  1737 => x"6e7e6b97",
  1738 => x"c880c148",
  1739 => x"98c758a6",
  1740 => x"7058a6cc",
  1741 => x"d2c37b97",
  1742 => x"87edfd87",
  1743 => x"87c28ef0",
  1744 => x"4c264d26",
  1745 => x"4f264b26",
  1746 => x"5c5b5e0e",
  1747 => x"86f40e5d",
  1748 => x"6d974d71",
  1749 => x"4ca5c17e",
  1750 => x"c8486c97",
  1751 => x"486e58a6",
  1752 => x"05a866c4",
  1753 => x"48ff87c5",
  1754 => x"fd87e6c0",
  1755 => x"a5c287c3",
  1756 => x"4b6c9749",
  1757 => x"974ba371",
  1758 => x"6c974b6b",
  1759 => x"c1486e7e",
  1760 => x"58a6c880",
  1761 => x"a6cc98c7",
  1762 => x"7c977058",
  1763 => x"7387dafc",
  1764 => x"fe8ef448",
  1765 => x"5e0e87ea",
  1766 => x"f40e5c5b",
  1767 => x"d84c7186",
  1768 => x"ffc34a66",
  1769 => x"4ba4c29a",
  1770 => x"73496c97",
  1771 => x"517249a1",
  1772 => x"6e7e6c97",
  1773 => x"c880c148",
  1774 => x"98c758a6",
  1775 => x"7058a6cc",
  1776 => x"fd8ef454",
  1777 => x"f01e87fc",
  1778 => x"7e699786",
  1779 => x"974aa1c1",
  1780 => x"a6c8486a",
  1781 => x"c4486e58",
  1782 => x"04a8b766",
  1783 => x"699787d3",
  1784 => x"486a977e",
  1785 => x"6e58a6c8",
  1786 => x"8866c448",
  1787 => x"d658a6cc",
  1788 => x"6e7e1187",
  1789 => x"a680c848",
  1790 => x"cc481258",
  1791 => x"66c458a6",
  1792 => x"8866c848",
  1793 => x"f058a6d0",
  1794 => x"1e4f268e",
  1795 => x"86f41e73",
  1796 => x"e087defa",
  1797 => x"c0494bbf",
  1798 => x"0299c0e0",
  1799 => x"1e7387cb",
  1800 => x"49cec6c3",
  1801 => x"c487effd",
  1802 => x"d0497386",
  1803 => x"c10299c0",
  1804 => x"c6c387c0",
  1805 => x"7ebf97d8",
  1806 => x"97d9c6c3",
  1807 => x"a6c848bf",
  1808 => x"c4486e58",
  1809 => x"c002a866",
  1810 => x"c6c387e8",
  1811 => x"49bf97d8",
  1812 => x"81dac6c3",
  1813 => x"08e04811",
  1814 => x"d8c6c378",
  1815 => x"6e7ebf97",
  1816 => x"c880c148",
  1817 => x"98c758a6",
  1818 => x"c358a6cc",
  1819 => x"c848d8c6",
  1820 => x"bfe45066",
  1821 => x"e0c0494b",
  1822 => x"cb0299c0",
  1823 => x"c31e7387",
  1824 => x"fc49e2c6",
  1825 => x"86c487d0",
  1826 => x"c0d04973",
  1827 => x"c0c10299",
  1828 => x"ecc6c387",
  1829 => x"c37ebf97",
  1830 => x"bf97edc6",
  1831 => x"58a6c848",
  1832 => x"66c4486e",
  1833 => x"e8c002a8",
  1834 => x"ecc6c387",
  1835 => x"c349bf97",
  1836 => x"1181eec6",
  1837 => x"7808e448",
  1838 => x"97ecc6c3",
  1839 => x"486e7ebf",
  1840 => x"a6c880c1",
  1841 => x"cc98c758",
  1842 => x"c6c358a6",
  1843 => x"66c848ec",
  1844 => x"87cbf750",
  1845 => x"d0f77e70",
  1846 => x"f98ef487",
  1847 => x"c31e87e6",
  1848 => x"f749cec6",
  1849 => x"c6c387d3",
  1850 => x"ccf749e2",
  1851 => x"cbf0c187",
  1852 => x"87dff649",
  1853 => x"2687c8c4",
  1854 => x"d0ff1e4f",
  1855 => x"78e1c848",
  1856 => x"c548d4ff",
  1857 => x"0266c478",
  1858 => x"e0c387c3",
  1859 => x"0266c878",
  1860 => x"d4ff87c6",
  1861 => x"78f0c348",
  1862 => x"7148d4ff",
  1863 => x"48d0ff78",
  1864 => x"c078e1c8",
  1865 => x"4f2678e0",
  1866 => x"5c5b5e0e",
  1867 => x"c34c710e",
  1868 => x"f849cec6",
  1869 => x"4a7087d2",
  1870 => x"04aab7c0",
  1871 => x"c387e3c2",
  1872 => x"c905aae0",
  1873 => x"f2f7c187",
  1874 => x"c278c148",
  1875 => x"f0c387d4",
  1876 => x"87c905aa",
  1877 => x"48eef7c1",
  1878 => x"f5c178c1",
  1879 => x"f2f7c187",
  1880 => x"87c702bf",
  1881 => x"c0c24b72",
  1882 => x"7287c2b3",
  1883 => x"059c744b",
  1884 => x"f7c187d1",
  1885 => x"c11ebfee",
  1886 => x"1ebff2f7",
  1887 => x"f8fd4972",
  1888 => x"c186c887",
  1889 => x"02bfeef7",
  1890 => x"7387e0c0",
  1891 => x"29b7c449",
  1892 => x"cef9c191",
  1893 => x"cf4a7381",
  1894 => x"c192c29a",
  1895 => x"70307248",
  1896 => x"72baff4a",
  1897 => x"70986948",
  1898 => x"7387db79",
  1899 => x"29b7c449",
  1900 => x"cef9c191",
  1901 => x"cf4a7381",
  1902 => x"c392c29a",
  1903 => x"70307248",
  1904 => x"b069484a",
  1905 => x"f7c17970",
  1906 => x"78c048f2",
  1907 => x"48eef7c1",
  1908 => x"c6c378c0",
  1909 => x"eff549ce",
  1910 => x"c04a7087",
  1911 => x"fd03aab7",
  1912 => x"48c087dd",
  1913 => x"4d2687c2",
  1914 => x"4b264c26",
  1915 => x"00004f26",
  1916 => x"00000000",
  1917 => x"711e0000",
  1918 => x"ebfc494a",
  1919 => x"1e4f2687",
  1920 => x"49724ac0",
  1921 => x"f9c191c4",
  1922 => x"79c081ce",
  1923 => x"b7d082c1",
  1924 => x"87ee04aa",
  1925 => x"5e0e4f26",
  1926 => x"0e5d5c5b",
  1927 => x"d0f24d71",
  1928 => x"c44a7587",
  1929 => x"c1922ab7",
  1930 => x"7582cef9",
  1931 => x"c29ccf4c",
  1932 => x"4b496a94",
  1933 => x"9bc32b74",
  1934 => x"307448c2",
  1935 => x"bcff4c70",
  1936 => x"98714874",
  1937 => x"e0f17a70",
  1938 => x"fe487387",
  1939 => x"000087d8",
  1940 => x"00000000",
  1941 => x"00000000",
  1942 => x"00000000",
  1943 => x"00000000",
  1944 => x"00000000",
  1945 => x"00000000",
  1946 => x"00000000",
  1947 => x"00000000",
  1948 => x"00000000",
  1949 => x"00000000",
  1950 => x"00000000",
  1951 => x"00000000",
  1952 => x"00000000",
  1953 => x"00000000",
  1954 => x"00000000",
  1955 => x"731e0000",
  1956 => x"c34b711e",
  1957 => x"f249e2c6",
  1958 => x"497087ee",
  1959 => x"49f0c11e",
  1960 => x"c487cbc8",
  1961 => x"e2c6c386",
  1962 => x"87dcf249",
  1963 => x"d4ff4970",
  1964 => x"c3787148",
  1965 => x"f249e2c6",
  1966 => x"497087ce",
  1967 => x"7148d4ff",
  1968 => x"05abc478",
  1969 => x"c6c387ce",
  1970 => x"fbf149e2",
  1971 => x"ff497087",
  1972 => x"787148d4",
  1973 => x"c048d0ff",
  1974 => x"87c478e0",
  1975 => x"4c264d26",
  1976 => x"4f264b26",
  1977 => x"5c5b5e0e",
  1978 => x"4a710e5d",
  1979 => x"87c6029a",
  1980 => x"48ffc1c2",
  1981 => x"c1c278c0",
  1982 => x"c105bfff",
  1983 => x"c6c387c6",
  1984 => x"c3f149e2",
  1985 => x"a8b7c087",
  1986 => x"c387cd04",
  1987 => x"f049e2c6",
  1988 => x"b7c087f6",
  1989 => x"87f303a8",
  1990 => x"bfffc1c2",
  1991 => x"ffc1c249",
  1992 => x"78a1c148",
  1993 => x"81cfc2c2",
  1994 => x"c2c24811",
  1995 => x"c2c258c7",
  1996 => x"78c048c7",
  1997 => x"c049f2c0",
  1998 => x"7087deec",
  1999 => x"fac6c349",
  2000 => x"87f8c459",
  2001 => x"bfc7c2c2",
  2002 => x"87f2c102",
  2003 => x"49e2c6c3",
  2004 => x"c087f5ef",
  2005 => x"cd04a8b7",
  2006 => x"c7c2c287",
  2007 => x"88c148bf",
  2008 => x"58cbc2c2",
  2009 => x"c6c387db",
  2010 => x"c049bff6",
  2011 => x"7087f6eb",
  2012 => x"87cd0298",
  2013 => x"49e2c6c3",
  2014 => x"c287feec",
  2015 => x"c048ffc1",
  2016 => x"c3c2c278",
  2017 => x"f3c305bf",
  2018 => x"c7c2c287",
  2019 => x"ebc305bf",
  2020 => x"ffc1c287",
  2021 => x"c1c249bf",
  2022 => x"a1c148ff",
  2023 => x"cfc2c278",
  2024 => x"494b1181",
  2025 => x"0299c0c2",
  2026 => x"7387ccc0",
  2027 => x"98ffc148",
  2028 => x"58cbc2c2",
  2029 => x"c287c5c3",
  2030 => x"c25bc7c2",
  2031 => x"c2c287fe",
  2032 => x"c102bfc3",
  2033 => x"c6c387db",
  2034 => x"c049bff6",
  2035 => x"7087d6ea",
  2036 => x"e7c20298",
  2037 => x"ffc1c287",
  2038 => x"c1c249bf",
  2039 => x"a1c148ff",
  2040 => x"cfc2c278",
  2041 => x"49699781",
  2042 => x"e2c6c31e",
  2043 => x"87e0eb49",
  2044 => x"c2c286c4",
  2045 => x"c149bfc3",
  2046 => x"c7c2c289",
  2047 => x"c7c2c259",
  2048 => x"7178c148",
  2049 => x"c6c00299",
  2050 => x"4cf2c087",
  2051 => x"d787c3c0",
  2052 => x"49744cdc",
  2053 => x"87c1e9c0",
  2054 => x"c6c34970",
  2055 => x"dbc159fa",
  2056 => x"e2c6c387",
  2057 => x"87deee49",
  2058 => x"029b4b70",
  2059 => x"c287eec0",
  2060 => x"b7bfcbc2",
  2061 => x"e4c003ab",
  2062 => x"f6c6c387",
  2063 => x"e8c049bf",
  2064 => x"987087e3",
  2065 => x"87f4c002",
  2066 => x"c2c248c7",
  2067 => x"c288bfcb",
  2068 => x"c358cfc2",
  2069 => x"e949e2c6",
  2070 => x"dfc087df",
  2071 => x"49dcd787",
  2072 => x"87f5e7c0",
  2073 => x"c6c34970",
  2074 => x"c2c259fa",
  2075 => x"b74abfcb",
  2076 => x"c7c004ab",
  2077 => x"d5f84987",
  2078 => x"87e5fe87",
  2079 => x"0087ddf9",
  2080 => x"00000000",
  2081 => x"00000000",
  2082 => x"04000000",
  2083 => x"01000000",
  2084 => x"f30882ff",
  2085 => x"f364f3c8",
  2086 => x"8101f250",
  2087 => x"1e00f401",
  2088 => x"c848d0ff",
  2089 => x"487178e1",
  2090 => x"7808d4ff",
  2091 => x"ff1e4f26",
  2092 => x"e1c848d0",
  2093 => x"ff487178",
  2094 => x"c47808d4",
  2095 => x"d4ff4866",
  2096 => x"4f267808",
  2097 => x"c44a711e",
  2098 => x"721e4966",
  2099 => x"87deff49",
  2100 => x"c048d0ff",
  2101 => x"262678e0",
  2102 => x"1e731e4f",
  2103 => x"66c84b71",
  2104 => x"4a731e49",
  2105 => x"49a2e0c1",
  2106 => x"2687d9ff",
  2107 => x"4d2687c4",
  2108 => x"4b264c26",
  2109 => x"ff1e4f26",
  2110 => x"ffc34ad4",
  2111 => x"48d0ff7a",
  2112 => x"de78e1c8",
  2113 => x"fac6c37a",
  2114 => x"48497abf",
  2115 => x"7a7028c8",
  2116 => x"28d04871",
  2117 => x"48717a70",
  2118 => x"7a7028d8",
  2119 => x"bffec6c3",
  2120 => x"c848497a",
  2121 => x"717a7028",
  2122 => x"7028d048",
  2123 => x"d848717a",
  2124 => x"ff7a7028",
  2125 => x"e0c048d0",
  2126 => x"1e4f2678",
  2127 => x"4a711e73",
  2128 => x"bffac6c3",
  2129 => x"c02b724b",
  2130 => x"ce04aae0",
  2131 => x"c0497287",
  2132 => x"c6c389e0",
  2133 => x"714bbffe",
  2134 => x"c087cf2b",
  2135 => x"897249e0",
  2136 => x"bffec6c3",
  2137 => x"70307148",
  2138 => x"66c8b349",
  2139 => x"c448739b",
  2140 => x"264d2687",
  2141 => x"264b264c",
  2142 => x"5b5e0e4f",
  2143 => x"ec0e5d5c",
  2144 => x"c34b7186",
  2145 => x"7ebffac6",
  2146 => x"c02c734c",
  2147 => x"c004abe0",
  2148 => x"a6c487e0",
  2149 => x"7378c048",
  2150 => x"89e0c049",
  2151 => x"e4c04a71",
  2152 => x"30724866",
  2153 => x"c358a6cc",
  2154 => x"4dbffec6",
  2155 => x"c02c714c",
  2156 => x"497387e4",
  2157 => x"4866e4c0",
  2158 => x"a6c83071",
  2159 => x"49e0c058",
  2160 => x"e4c08973",
  2161 => x"28714866",
  2162 => x"c358a6cc",
  2163 => x"4dbffec6",
  2164 => x"70307148",
  2165 => x"e4c0b449",
  2166 => x"84c19c66",
  2167 => x"ac66e8c0",
  2168 => x"c087c204",
  2169 => x"abe0c04c",
  2170 => x"cc87d304",
  2171 => x"78c048a6",
  2172 => x"e0c04973",
  2173 => x"71487489",
  2174 => x"58a6d430",
  2175 => x"497387d5",
  2176 => x"30714874",
  2177 => x"c058a6d0",
  2178 => x"897349e0",
  2179 => x"28714874",
  2180 => x"c458a6d4",
  2181 => x"baff4a66",
  2182 => x"66c89a6e",
  2183 => x"75b9ff49",
  2184 => x"cc487299",
  2185 => x"c6c3b066",
  2186 => x"487158fe",
  2187 => x"c3b066d0",
  2188 => x"fb58c2c7",
  2189 => x"8eec87c0",
  2190 => x"1e87f6fc",
  2191 => x"c848d0ff",
  2192 => x"487178c9",
  2193 => x"7808d4ff",
  2194 => x"711e4f26",
  2195 => x"87eb494a",
  2196 => x"c848d0ff",
  2197 => x"1e4f2678",
  2198 => x"4b711e73",
  2199 => x"bfcec7c3",
  2200 => x"c287c302",
  2201 => x"d0ff87eb",
  2202 => x"78c9c848",
  2203 => x"e0c04973",
  2204 => x"48d4ffb1",
  2205 => x"c7c37871",
  2206 => x"78c048c2",
  2207 => x"c50266c8",
  2208 => x"49ffc387",
  2209 => x"49c087c2",
  2210 => x"59cac7c3",
  2211 => x"c60266cc",
  2212 => x"d5d5c587",
  2213 => x"cf87c44a",
  2214 => x"c34affff",
  2215 => x"c35acec7",
  2216 => x"c148cec7",
  2217 => x"2687c478",
  2218 => x"264c264d",
  2219 => x"0e4f264b",
  2220 => x"5d5c5b5e",
  2221 => x"c34a710e",
  2222 => x"4cbfcac7",
  2223 => x"cb029a72",
  2224 => x"91c84987",
  2225 => x"4bcdc9c2",
  2226 => x"87c48371",
  2227 => x"4bcdcdc2",
  2228 => x"49134dc0",
  2229 => x"c7c39974",
  2230 => x"ffb9bfc6",
  2231 => x"787148d4",
  2232 => x"852cb7c1",
  2233 => x"04adb7c8",
  2234 => x"c7c387e8",
  2235 => x"c848bfc2",
  2236 => x"c6c7c380",
  2237 => x"87effe58",
  2238 => x"711e731e",
  2239 => x"9a4a134b",
  2240 => x"7287cb02",
  2241 => x"87e7fe49",
  2242 => x"059a4a13",
  2243 => x"dafe87f5",
  2244 => x"c7c31e87",
  2245 => x"c349bfc2",
  2246 => x"c148c2c7",
  2247 => x"c0c478a1",
  2248 => x"db03a9b7",
  2249 => x"48d4ff87",
  2250 => x"bfc6c7c3",
  2251 => x"c2c7c378",
  2252 => x"c7c349bf",
  2253 => x"a1c148c2",
  2254 => x"b7c0c478",
  2255 => x"87e504a9",
  2256 => x"c848d0ff",
  2257 => x"cec7c378",
  2258 => x"2678c048",
  2259 => x"0000004f",
  2260 => x"00000000",
  2261 => x"00000000",
  2262 => x"00005f5f",
  2263 => x"03030000",
  2264 => x"00030300",
  2265 => x"7f7f1400",
  2266 => x"147f7f14",
  2267 => x"2e240000",
  2268 => x"123a6b6b",
  2269 => x"366a4c00",
  2270 => x"32566c18",
  2271 => x"4f7e3000",
  2272 => x"683a7759",
  2273 => x"04000040",
  2274 => x"00000307",
  2275 => x"1c000000",
  2276 => x"0041633e",
  2277 => x"41000000",
  2278 => x"001c3e63",
  2279 => x"3e2a0800",
  2280 => x"2a3e1c1c",
  2281 => x"08080008",
  2282 => x"08083e3e",
  2283 => x"80000000",
  2284 => x"000060e0",
  2285 => x"08080000",
  2286 => x"08080808",
  2287 => x"00000000",
  2288 => x"00006060",
  2289 => x"30604000",
  2290 => x"03060c18",
  2291 => x"7f3e0001",
  2292 => x"3e7f4d59",
  2293 => x"06040000",
  2294 => x"00007f7f",
  2295 => x"63420000",
  2296 => x"464f5971",
  2297 => x"63220000",
  2298 => x"367f4949",
  2299 => x"161c1800",
  2300 => x"107f7f13",
  2301 => x"67270000",
  2302 => x"397d4545",
  2303 => x"7e3c0000",
  2304 => x"3079494b",
  2305 => x"01010000",
  2306 => x"070f7971",
  2307 => x"7f360000",
  2308 => x"367f4949",
  2309 => x"4f060000",
  2310 => x"1e3f6949",
  2311 => x"00000000",
  2312 => x"00006666",
  2313 => x"80000000",
  2314 => x"000066e6",
  2315 => x"08080000",
  2316 => x"22221414",
  2317 => x"14140000",
  2318 => x"14141414",
  2319 => x"22220000",
  2320 => x"08081414",
  2321 => x"03020000",
  2322 => x"060f5951",
  2323 => x"417f3e00",
  2324 => x"1e1f555d",
  2325 => x"7f7e0000",
  2326 => x"7e7f0909",
  2327 => x"7f7f0000",
  2328 => x"367f4949",
  2329 => x"3e1c0000",
  2330 => x"41414163",
  2331 => x"7f7f0000",
  2332 => x"1c3e6341",
  2333 => x"7f7f0000",
  2334 => x"41414949",
  2335 => x"7f7f0000",
  2336 => x"01010909",
  2337 => x"7f3e0000",
  2338 => x"7a7b4941",
  2339 => x"7f7f0000",
  2340 => x"7f7f0808",
  2341 => x"41000000",
  2342 => x"00417f7f",
  2343 => x"60200000",
  2344 => x"3f7f4040",
  2345 => x"087f7f00",
  2346 => x"4163361c",
  2347 => x"7f7f0000",
  2348 => x"40404040",
  2349 => x"067f7f00",
  2350 => x"7f7f060c",
  2351 => x"067f7f00",
  2352 => x"7f7f180c",
  2353 => x"7f3e0000",
  2354 => x"3e7f4141",
  2355 => x"7f7f0000",
  2356 => x"060f0909",
  2357 => x"417f3e00",
  2358 => x"407e7f61",
  2359 => x"7f7f0000",
  2360 => x"667f1909",
  2361 => x"6f260000",
  2362 => x"327b594d",
  2363 => x"01010000",
  2364 => x"01017f7f",
  2365 => x"7f3f0000",
  2366 => x"3f7f4040",
  2367 => x"3f0f0000",
  2368 => x"0f3f7070",
  2369 => x"307f7f00",
  2370 => x"7f7f3018",
  2371 => x"36634100",
  2372 => x"63361c1c",
  2373 => x"06030141",
  2374 => x"03067c7c",
  2375 => x"59716101",
  2376 => x"4143474d",
  2377 => x"7f000000",
  2378 => x"0041417f",
  2379 => x"06030100",
  2380 => x"6030180c",
  2381 => x"41000040",
  2382 => x"007f7f41",
  2383 => x"060c0800",
  2384 => x"080c0603",
  2385 => x"80808000",
  2386 => x"80808080",
  2387 => x"00000000",
  2388 => x"00040703",
  2389 => x"74200000",
  2390 => x"787c5454",
  2391 => x"7f7f0000",
  2392 => x"387c4444",
  2393 => x"7c380000",
  2394 => x"00444444",
  2395 => x"7c380000",
  2396 => x"7f7f4444",
  2397 => x"7c380000",
  2398 => x"185c5454",
  2399 => x"7e040000",
  2400 => x"0005057f",
  2401 => x"bc180000",
  2402 => x"7cfca4a4",
  2403 => x"7f7f0000",
  2404 => x"787c0404",
  2405 => x"00000000",
  2406 => x"00407d3d",
  2407 => x"80800000",
  2408 => x"007dfd80",
  2409 => x"7f7f0000",
  2410 => x"446c3810",
  2411 => x"00000000",
  2412 => x"00407f3f",
  2413 => x"0c7c7c00",
  2414 => x"787c0c18",
  2415 => x"7c7c0000",
  2416 => x"787c0404",
  2417 => x"7c380000",
  2418 => x"387c4444",
  2419 => x"fcfc0000",
  2420 => x"183c2424",
  2421 => x"3c180000",
  2422 => x"fcfc2424",
  2423 => x"7c7c0000",
  2424 => x"080c0404",
  2425 => x"5c480000",
  2426 => x"20745454",
  2427 => x"3f040000",
  2428 => x"0044447f",
  2429 => x"7c3c0000",
  2430 => x"7c7c4040",
  2431 => x"3c1c0000",
  2432 => x"1c3c6060",
  2433 => x"607c3c00",
  2434 => x"3c7c6030",
  2435 => x"386c4400",
  2436 => x"446c3810",
  2437 => x"bc1c0000",
  2438 => x"1c3c60e0",
  2439 => x"64440000",
  2440 => x"444c5c74",
  2441 => x"08080000",
  2442 => x"4141773e",
  2443 => x"00000000",
  2444 => x"00007f7f",
  2445 => x"41410000",
  2446 => x"08083e77",
  2447 => x"01010200",
  2448 => x"01020203",
  2449 => x"7f7f7f00",
  2450 => x"7f7f7f7f",
  2451 => x"1c080800",
  2452 => x"7f3e3e1c",
  2453 => x"3e7f7f7f",
  2454 => x"081c1c3e",
  2455 => x"18100008",
  2456 => x"10187c7c",
  2457 => x"30100000",
  2458 => x"10307c7c",
  2459 => x"60301000",
  2460 => x"061e7860",
  2461 => x"3c664200",
  2462 => x"42663c18",
  2463 => x"6a387800",
  2464 => x"386cc6c2",
  2465 => x"00006000",
  2466 => x"60000060",
  2467 => x"5b5e0e00",
  2468 => x"1e0e5d5c",
  2469 => x"c7c34c71",
  2470 => x"c04dbfdf",
  2471 => x"741ec04b",
  2472 => x"87c702ab",
  2473 => x"c048a6c4",
  2474 => x"c487c578",
  2475 => x"78c148a6",
  2476 => x"731e66c4",
  2477 => x"87dfee49",
  2478 => x"e0c086c8",
  2479 => x"87efef49",
  2480 => x"6a4aa5c4",
  2481 => x"87f0f049",
  2482 => x"cb87c6f1",
  2483 => x"c883c185",
  2484 => x"ff04abb7",
  2485 => x"262687c7",
  2486 => x"264c264d",
  2487 => x"1e4f264b",
  2488 => x"c7c34a71",
  2489 => x"c7c35ae3",
  2490 => x"78c748e3",
  2491 => x"87ddfe49",
  2492 => x"731e4f26",
  2493 => x"c04a711e",
  2494 => x"d303aab7",
  2495 => x"d1e9c287",
  2496 => x"87c405bf",
  2497 => x"87c24bc1",
  2498 => x"e9c24bc0",
  2499 => x"87c45bd5",
  2500 => x"5ad5e9c2",
  2501 => x"bfd1e9c2",
  2502 => x"c19ac14a",
  2503 => x"ec49a2c0",
  2504 => x"48fc87e8",
  2505 => x"bfd1e9c2",
  2506 => x"87effe78",
  2507 => x"c44a711e",
  2508 => x"49721e66",
  2509 => x"2687e2e6",
  2510 => x"c21e4f26",
  2511 => x"49bfd1e9",
  2512 => x"87f2daff",
  2513 => x"48d7c7c3",
  2514 => x"c378bfe8",
  2515 => x"ec48d3c7",
  2516 => x"c7c378bf",
  2517 => x"494abfd7",
  2518 => x"c899ffc3",
  2519 => x"48722ab7",
  2520 => x"c7c3b071",
  2521 => x"4f2658df",
  2522 => x"5c5b5e0e",
  2523 => x"4b710e5d",
  2524 => x"c387c7ff",
  2525 => x"c048d2c7",
  2526 => x"ff497350",
  2527 => x"7087d7da",
  2528 => x"9cc24c49",
  2529 => x"cb49eecb",
  2530 => x"497087cf",
  2531 => x"d2c7c34d",
  2532 => x"c105bf97",
  2533 => x"66d087e4",
  2534 => x"dbc7c349",
  2535 => x"d70599bf",
  2536 => x"4966d487",
  2537 => x"bfd3c7c3",
  2538 => x"87cc0599",
  2539 => x"d9ff4973",
  2540 => x"987087e4",
  2541 => x"87c2c102",
  2542 => x"fdfd4cc1",
  2543 => x"ca497587",
  2544 => x"987087e3",
  2545 => x"c387c602",
  2546 => x"c148d2c7",
  2547 => x"d2c7c350",
  2548 => x"c005bf97",
  2549 => x"c7c387e4",
  2550 => x"d049bfdb",
  2551 => x"ff059966",
  2552 => x"c7c387d6",
  2553 => x"d449bfd3",
  2554 => x"ff059966",
  2555 => x"497387ca",
  2556 => x"87e2d8ff",
  2557 => x"fe059870",
  2558 => x"487487fe",
  2559 => x"0e87d8fb",
  2560 => x"5d5c5b5e",
  2561 => x"c086f40e",
  2562 => x"bfec4c4d",
  2563 => x"48a6c47e",
  2564 => x"bfdfc7c3",
  2565 => x"c01ec178",
  2566 => x"fd49c71e",
  2567 => x"86c887ca",
  2568 => x"ce029870",
  2569 => x"fb49ff87",
  2570 => x"dac187c8",
  2571 => x"e5d7ff49",
  2572 => x"c34dc187",
  2573 => x"bf97d2c7",
  2574 => x"d087c302",
  2575 => x"c7c387c5",
  2576 => x"c24bbfd7",
  2577 => x"05bfd1e9",
  2578 => x"c387ebc0",
  2579 => x"d7ff49fd",
  2580 => x"fac387c4",
  2581 => x"fdd6ff49",
  2582 => x"c3497387",
  2583 => x"1e7199ff",
  2584 => x"c7fb49c0",
  2585 => x"c8497387",
  2586 => x"1e7129b7",
  2587 => x"fbfa49c1",
  2588 => x"c686c887",
  2589 => x"c7c387c1",
  2590 => x"9b4bbfdb",
  2591 => x"c287dd02",
  2592 => x"49bfcde9",
  2593 => x"7087dec7",
  2594 => x"87c40598",
  2595 => x"87d24bc0",
  2596 => x"c749e0c2",
  2597 => x"e9c287c3",
  2598 => x"87c658d1",
  2599 => x"48cde9c2",
  2600 => x"497378c0",
  2601 => x"ce0599c2",
  2602 => x"49ebc387",
  2603 => x"87e6d5ff",
  2604 => x"99c24970",
  2605 => x"fb87c202",
  2606 => x"c149734c",
  2607 => x"87ce0599",
  2608 => x"ff49f4c3",
  2609 => x"7087cfd5",
  2610 => x"0299c249",
  2611 => x"4cfa87c2",
  2612 => x"99c84973",
  2613 => x"c387ce05",
  2614 => x"d4ff49f5",
  2615 => x"497087f8",
  2616 => x"d50299c2",
  2617 => x"e3c7c387",
  2618 => x"87ca02bf",
  2619 => x"c388c148",
  2620 => x"c058e7c7",
  2621 => x"4cff87c2",
  2622 => x"49734dc1",
  2623 => x"ce0599c4",
  2624 => x"49f2c387",
  2625 => x"87ced4ff",
  2626 => x"99c24970",
  2627 => x"c387dc02",
  2628 => x"7ebfe3c7",
  2629 => x"a8b7c748",
  2630 => x"87cbc003",
  2631 => x"80c1486e",
  2632 => x"58e7c7c3",
  2633 => x"fe87c2c0",
  2634 => x"c34dc14c",
  2635 => x"d3ff49fd",
  2636 => x"497087e4",
  2637 => x"c00299c2",
  2638 => x"c7c387d5",
  2639 => x"c002bfe3",
  2640 => x"c7c387c9",
  2641 => x"78c048e3",
  2642 => x"fd87c2c0",
  2643 => x"c34dc14c",
  2644 => x"d3ff49fa",
  2645 => x"497087c0",
  2646 => x"c00299c2",
  2647 => x"c7c387d9",
  2648 => x"c748bfe3",
  2649 => x"c003a8b7",
  2650 => x"c7c387c9",
  2651 => x"78c748e3",
  2652 => x"fc87c2c0",
  2653 => x"c04dc14c",
  2654 => x"c003acb7",
  2655 => x"66c487d1",
  2656 => x"82d8c14a",
  2657 => x"c6c0026a",
  2658 => x"744b6a87",
  2659 => x"c00f7349",
  2660 => x"1ef0c31e",
  2661 => x"f749dac1",
  2662 => x"86c887ce",
  2663 => x"c0029870",
  2664 => x"a6c887e2",
  2665 => x"e3c7c348",
  2666 => x"66c878bf",
  2667 => x"c491cb49",
  2668 => x"80714866",
  2669 => x"bf6e7e70",
  2670 => x"87c8c002",
  2671 => x"c84bbf6e",
  2672 => x"0f734966",
  2673 => x"c0029d75",
  2674 => x"c7c387c8",
  2675 => x"f249bfe3",
  2676 => x"e9c287fb",
  2677 => x"c002bfd5",
  2678 => x"c24987dd",
  2679 => x"987087c7",
  2680 => x"87d3c002",
  2681 => x"bfe3c7c3",
  2682 => x"87e1f249",
  2683 => x"c1f449c0",
  2684 => x"d5e9c287",
  2685 => x"f478c048",
  2686 => x"87dbf38e",
  2687 => x"5c5b5e0e",
  2688 => x"711e0e5d",
  2689 => x"dfc7c34c",
  2690 => x"cdc149bf",
  2691 => x"d1c14da1",
  2692 => x"747e6981",
  2693 => x"87cf029c",
  2694 => x"744ba5c4",
  2695 => x"dfc7c37b",
  2696 => x"faf249bf",
  2697 => x"747b6e87",
  2698 => x"87c4059c",
  2699 => x"87c24bc0",
  2700 => x"49734bc1",
  2701 => x"d487fbf2",
  2702 => x"87c70266",
  2703 => x"7087da49",
  2704 => x"c087c24a",
  2705 => x"d9e9c24a",
  2706 => x"caf2265a",
  2707 => x"00000087",
  2708 => x"00000000",
  2709 => x"00000000",
  2710 => x"4a711e00",
  2711 => x"49bfc8ff",
  2712 => x"2648a172",
  2713 => x"c8ff1e4f",
  2714 => x"c0fe89bf",
  2715 => x"c0c0c0c0",
  2716 => x"87c401a9",
  2717 => x"87c24ac0",
  2718 => x"48724ac1",
  2719 => x"5e0e4f26",
  2720 => x"0e5d5c5b",
  2721 => x"d4ff4b71",
  2722 => x"4866d04c",
  2723 => x"49d678c0",
  2724 => x"87cbd8ff",
  2725 => x"6c7cffc3",
  2726 => x"99ffc349",
  2727 => x"c3494d71",
  2728 => x"e0c199f0",
  2729 => x"87cb05a9",
  2730 => x"6c7cffc3",
  2731 => x"d098c348",
  2732 => x"c3780866",
  2733 => x"4a6c7cff",
  2734 => x"c331c849",
  2735 => x"4a6c7cff",
  2736 => x"4972b271",
  2737 => x"ffc331c8",
  2738 => x"714a6c7c",
  2739 => x"c84972b2",
  2740 => x"7cffc331",
  2741 => x"b2714a6c",
  2742 => x"c048d0ff",
  2743 => x"9b7378e0",
  2744 => x"7287c202",
  2745 => x"2648757b",
  2746 => x"264c264d",
  2747 => x"1e4f264b",
  2748 => x"5e0e4f26",
  2749 => x"f80e5c5b",
  2750 => x"c81e7686",
  2751 => x"fdfd49a6",
  2752 => x"7086c487",
  2753 => x"c2486e4b",
  2754 => x"f0c203a8",
  2755 => x"c34a7387",
  2756 => x"d0c19af0",
  2757 => x"87c702aa",
  2758 => x"05aae0c1",
  2759 => x"7387dec2",
  2760 => x"0299c849",
  2761 => x"c6ff87c3",
  2762 => x"c34c7387",
  2763 => x"05acc29c",
  2764 => x"c487c2c1",
  2765 => x"31c94966",
  2766 => x"66c41e71",
  2767 => x"c392d44a",
  2768 => x"7249e7c7",
  2769 => x"d7fafd81",
  2770 => x"ff49d887",
  2771 => x"c887d0d5",
  2772 => x"f5c21ec0",
  2773 => x"d6fd49de",
  2774 => x"d0ff87d2",
  2775 => x"78e0c048",
  2776 => x"1edef5c2",
  2777 => x"d44a66cc",
  2778 => x"e7c7c392",
  2779 => x"fd817249",
  2780 => x"cc87def8",
  2781 => x"05acc186",
  2782 => x"c487c2c1",
  2783 => x"31c94966",
  2784 => x"66c41e71",
  2785 => x"c392d44a",
  2786 => x"7249e7c7",
  2787 => x"cff9fd81",
  2788 => x"def5c287",
  2789 => x"4a66c81e",
  2790 => x"c7c392d4",
  2791 => x"817249e7",
  2792 => x"87def6fd",
  2793 => x"d3ff49d7",
  2794 => x"c0c887f5",
  2795 => x"def5c21e",
  2796 => x"d0d4fd49",
  2797 => x"ff86cc87",
  2798 => x"e0c048d0",
  2799 => x"fc8ef878",
  2800 => x"5e0e87e7",
  2801 => x"0e5d5c5b",
  2802 => x"ff4d711e",
  2803 => x"66d44cd4",
  2804 => x"b7c3487e",
  2805 => x"87c506a8",
  2806 => x"e2c148c0",
  2807 => x"fe497587",
  2808 => x"7587e3c7",
  2809 => x"4b66c41e",
  2810 => x"c7c393d4",
  2811 => x"497383e7",
  2812 => x"87f9f1fd",
  2813 => x"4b6b83c8",
  2814 => x"c848d0ff",
  2815 => x"7cdd78e1",
  2816 => x"ffc34973",
  2817 => x"737c7199",
  2818 => x"29b7c849",
  2819 => x"7199ffc3",
  2820 => x"d049737c",
  2821 => x"ffc329b7",
  2822 => x"737c7199",
  2823 => x"29b7d849",
  2824 => x"7cc07c71",
  2825 => x"7c7c7c7c",
  2826 => x"7c7c7c7c",
  2827 => x"c07c7c7c",
  2828 => x"66c478e0",
  2829 => x"ff49dc1e",
  2830 => x"c887c9d2",
  2831 => x"26487386",
  2832 => x"1e87e4fa",
  2833 => x"bff4f4c2",
  2834 => x"c2b9c149",
  2835 => x"ff59f8f4",
  2836 => x"ffc348d4",
  2837 => x"48d0ff78",
  2838 => x"ff78e1c8",
  2839 => x"78c148d4",
  2840 => x"787131c4",
  2841 => x"c048d0ff",
  2842 => x"4f2678e0",
  2843 => x"c5f2c21e",
  2844 => x"d4c2c31e",
  2845 => x"f4effd49",
  2846 => x"7086c487",
  2847 => x"87c30298",
  2848 => x"2687c0ff",
  2849 => x"4b35314f",
  2850 => x"20205a48",
  2851 => x"47464320",
  2852 => x"4a711e00",
  2853 => x"c349a2c4",
  2854 => x"6a48fac6",
  2855 => x"c1496978",
  2856 => x"f8f4c2b9",
  2857 => x"87dbfe59",
  2858 => x"87cad1ff",
  2859 => x"4f2648c1",
  2860 => x"c44a711e",
  2861 => x"c6c349a2",
  2862 => x"c27abffa",
  2863 => x"79bff4f4",
  2864 => x"711e4f26",
  2865 => x"c0029a4a",
  2866 => x"c31e87ec",
  2867 => x"fd49d4c2",
  2868 => x"c487daee",
  2869 => x"02987086",
  2870 => x"f5c287dc",
  2871 => x"c2c31ede",
  2872 => x"f1fd49d4",
  2873 => x"86c487dc",
  2874 => x"c9029870",
  2875 => x"def5c287",
  2876 => x"87ddfe49",
  2877 => x"48c087c2",
  2878 => x"711e4f26",
  2879 => x"c0029a4a",
  2880 => x"c31e87ee",
  2881 => x"fd49d4c2",
  2882 => x"c487e2ed",
  2883 => x"02987086",
  2884 => x"f5c287de",
  2885 => x"d7fe49de",
  2886 => x"def5c287",
  2887 => x"d4c2c31e",
  2888 => x"ecf1fd49",
  2889 => x"7086c487",
  2890 => x"87c40298",
  2891 => x"87c248c1",
  2892 => x"4f2648c0",
  2893 => x"00000000",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
