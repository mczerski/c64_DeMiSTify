library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom2 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"7178c148",
     1 => x"c6c00299",
     2 => x"4cf2c087",
     3 => x"d787c3c0",
     4 => x"49744cdc",
     5 => x"87c1e9c0",
     6 => x"c6c34970",
     7 => x"dbc159fa",
     8 => x"e2c6c387",
     9 => x"87deee49",
    10 => x"029b4b70",
    11 => x"c287eec0",
    12 => x"b7bfcbc2",
    13 => x"e4c003ab",
    14 => x"f6c6c387",
    15 => x"e8c049bf",
    16 => x"987087e3",
    17 => x"87f4c002",
    18 => x"c2c248c7",
    19 => x"c288bfcb",
    20 => x"c358cfc2",
    21 => x"e949e2c6",
    22 => x"dfc087df",
    23 => x"49dcd787",
    24 => x"87f5e7c0",
    25 => x"c6c34970",
    26 => x"c2c259fa",
    27 => x"b74abfcb",
    28 => x"c7c004ab",
    29 => x"d5f84987",
    30 => x"87e5fe87",
    31 => x"0087ddf9",
    32 => x"00000000",
    33 => x"00000000",
    34 => x"04000000",
    35 => x"01000000",
    36 => x"f30882ff",
    37 => x"f364f3c8",
    38 => x"8101f250",
    39 => x"1e00f401",
    40 => x"c848d0ff",
    41 => x"487178e1",
    42 => x"7808d4ff",
    43 => x"ff1e4f26",
    44 => x"e1c848d0",
    45 => x"ff487178",
    46 => x"c47808d4",
    47 => x"d4ff4866",
    48 => x"4f267808",
    49 => x"c44a711e",
    50 => x"721e4966",
    51 => x"87deff49",
    52 => x"c048d0ff",
    53 => x"262678e0",
    54 => x"1e731e4f",
    55 => x"66c84b71",
    56 => x"4a731e49",
    57 => x"49a2e0c1",
    58 => x"2687d9ff",
    59 => x"4d2687c4",
    60 => x"4b264c26",
    61 => x"ff1e4f26",
    62 => x"ffc34ad4",
    63 => x"48d0ff7a",
    64 => x"de78e1c8",
    65 => x"fac6c37a",
    66 => x"48497abf",
    67 => x"7a7028c8",
    68 => x"28d04871",
    69 => x"48717a70",
    70 => x"7a7028d8",
    71 => x"bffec6c3",
    72 => x"c848497a",
    73 => x"717a7028",
    74 => x"7028d048",
    75 => x"d848717a",
    76 => x"ff7a7028",
    77 => x"e0c048d0",
    78 => x"1e4f2678",
    79 => x"4a711e73",
    80 => x"bffac6c3",
    81 => x"c02b724b",
    82 => x"ce04aae0",
    83 => x"c0497287",
    84 => x"c6c389e0",
    85 => x"714bbffe",
    86 => x"c087cf2b",
    87 => x"897249e0",
    88 => x"bffec6c3",
    89 => x"70307148",
    90 => x"66c8b349",
    91 => x"c448739b",
    92 => x"264d2687",
    93 => x"264b264c",
    94 => x"5b5e0e4f",
    95 => x"ec0e5d5c",
    96 => x"c34b7186",
    97 => x"7ebffac6",
    98 => x"c02c734c",
    99 => x"c004abe0",
   100 => x"a6c487e0",
   101 => x"7378c048",
   102 => x"89e0c049",
   103 => x"e4c04a71",
   104 => x"30724866",
   105 => x"c358a6cc",
   106 => x"4dbffec6",
   107 => x"c02c714c",
   108 => x"497387e4",
   109 => x"4866e4c0",
   110 => x"a6c83071",
   111 => x"49e0c058",
   112 => x"e4c08973",
   113 => x"28714866",
   114 => x"c358a6cc",
   115 => x"4dbffec6",
   116 => x"70307148",
   117 => x"e4c0b449",
   118 => x"84c19c66",
   119 => x"ac66e8c0",
   120 => x"c087c204",
   121 => x"abe0c04c",
   122 => x"cc87d304",
   123 => x"78c048a6",
   124 => x"e0c04973",
   125 => x"71487489",
   126 => x"58a6d430",
   127 => x"497387d5",
   128 => x"30714874",
   129 => x"c058a6d0",
   130 => x"897349e0",
   131 => x"28714874",
   132 => x"c458a6d4",
   133 => x"baff4a66",
   134 => x"66c89a6e",
   135 => x"75b9ff49",
   136 => x"cc487299",
   137 => x"c6c3b066",
   138 => x"487158fe",
   139 => x"c3b066d0",
   140 => x"fb58c2c7",
   141 => x"8eec87c0",
   142 => x"1e87f6fc",
   143 => x"c848d0ff",
   144 => x"487178c9",
   145 => x"7808d4ff",
   146 => x"711e4f26",
   147 => x"87eb494a",
   148 => x"c848d0ff",
   149 => x"1e4f2678",
   150 => x"4b711e73",
   151 => x"bfcec7c3",
   152 => x"c287c302",
   153 => x"d0ff87eb",
   154 => x"78c9c848",
   155 => x"e0c04973",
   156 => x"48d4ffb1",
   157 => x"c7c37871",
   158 => x"78c048c2",
   159 => x"c50266c8",
   160 => x"49ffc387",
   161 => x"49c087c2",
   162 => x"59cac7c3",
   163 => x"c60266cc",
   164 => x"d5d5c587",
   165 => x"cf87c44a",
   166 => x"c34affff",
   167 => x"c35acec7",
   168 => x"c148cec7",
   169 => x"2687c478",
   170 => x"264c264d",
   171 => x"0e4f264b",
   172 => x"5d5c5b5e",
   173 => x"c34a710e",
   174 => x"4cbfcac7",
   175 => x"cb029a72",
   176 => x"91c84987",
   177 => x"4bcdc9c2",
   178 => x"87c48371",
   179 => x"4bcdcdc2",
   180 => x"49134dc0",
   181 => x"c7c39974",
   182 => x"ffb9bfc6",
   183 => x"787148d4",
   184 => x"852cb7c1",
   185 => x"04adb7c8",
   186 => x"c7c387e8",
   187 => x"c848bfc2",
   188 => x"c6c7c380",
   189 => x"87effe58",
   190 => x"711e731e",
   191 => x"9a4a134b",
   192 => x"7287cb02",
   193 => x"87e7fe49",
   194 => x"059a4a13",
   195 => x"dafe87f5",
   196 => x"c7c31e87",
   197 => x"c349bfc2",
   198 => x"c148c2c7",
   199 => x"c0c478a1",
   200 => x"db03a9b7",
   201 => x"48d4ff87",
   202 => x"bfc6c7c3",
   203 => x"c2c7c378",
   204 => x"c7c349bf",
   205 => x"a1c148c2",
   206 => x"b7c0c478",
   207 => x"87e504a9",
   208 => x"c848d0ff",
   209 => x"cec7c378",
   210 => x"2678c048",
   211 => x"0000004f",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00005f5f",
   215 => x"03030000",
   216 => x"00030300",
   217 => x"7f7f1400",
   218 => x"147f7f14",
   219 => x"2e240000",
   220 => x"123a6b6b",
   221 => x"366a4c00",
   222 => x"32566c18",
   223 => x"4f7e3000",
   224 => x"683a7759",
   225 => x"04000040",
   226 => x"00000307",
   227 => x"1c000000",
   228 => x"0041633e",
   229 => x"41000000",
   230 => x"001c3e63",
   231 => x"3e2a0800",
   232 => x"2a3e1c1c",
   233 => x"08080008",
   234 => x"08083e3e",
   235 => x"80000000",
   236 => x"000060e0",
   237 => x"08080000",
   238 => x"08080808",
   239 => x"00000000",
   240 => x"00006060",
   241 => x"30604000",
   242 => x"03060c18",
   243 => x"7f3e0001",
   244 => x"3e7f4d59",
   245 => x"06040000",
   246 => x"00007f7f",
   247 => x"63420000",
   248 => x"464f5971",
   249 => x"63220000",
   250 => x"367f4949",
   251 => x"161c1800",
   252 => x"107f7f13",
   253 => x"67270000",
   254 => x"397d4545",
   255 => x"7e3c0000",
   256 => x"3079494b",
   257 => x"01010000",
   258 => x"070f7971",
   259 => x"7f360000",
   260 => x"367f4949",
   261 => x"4f060000",
   262 => x"1e3f6949",
   263 => x"00000000",
   264 => x"00006666",
   265 => x"80000000",
   266 => x"000066e6",
   267 => x"08080000",
   268 => x"22221414",
   269 => x"14140000",
   270 => x"14141414",
   271 => x"22220000",
   272 => x"08081414",
   273 => x"03020000",
   274 => x"060f5951",
   275 => x"417f3e00",
   276 => x"1e1f555d",
   277 => x"7f7e0000",
   278 => x"7e7f0909",
   279 => x"7f7f0000",
   280 => x"367f4949",
   281 => x"3e1c0000",
   282 => x"41414163",
   283 => x"7f7f0000",
   284 => x"1c3e6341",
   285 => x"7f7f0000",
   286 => x"41414949",
   287 => x"7f7f0000",
   288 => x"01010909",
   289 => x"7f3e0000",
   290 => x"7a7b4941",
   291 => x"7f7f0000",
   292 => x"7f7f0808",
   293 => x"41000000",
   294 => x"00417f7f",
   295 => x"60200000",
   296 => x"3f7f4040",
   297 => x"087f7f00",
   298 => x"4163361c",
   299 => x"7f7f0000",
   300 => x"40404040",
   301 => x"067f7f00",
   302 => x"7f7f060c",
   303 => x"067f7f00",
   304 => x"7f7f180c",
   305 => x"7f3e0000",
   306 => x"3e7f4141",
   307 => x"7f7f0000",
   308 => x"060f0909",
   309 => x"417f3e00",
   310 => x"407e7f61",
   311 => x"7f7f0000",
   312 => x"667f1909",
   313 => x"6f260000",
   314 => x"327b594d",
   315 => x"01010000",
   316 => x"01017f7f",
   317 => x"7f3f0000",
   318 => x"3f7f4040",
   319 => x"3f0f0000",
   320 => x"0f3f7070",
   321 => x"307f7f00",
   322 => x"7f7f3018",
   323 => x"36634100",
   324 => x"63361c1c",
   325 => x"06030141",
   326 => x"03067c7c",
   327 => x"59716101",
   328 => x"4143474d",
   329 => x"7f000000",
   330 => x"0041417f",
   331 => x"06030100",
   332 => x"6030180c",
   333 => x"41000040",
   334 => x"007f7f41",
   335 => x"060c0800",
   336 => x"080c0603",
   337 => x"80808000",
   338 => x"80808080",
   339 => x"00000000",
   340 => x"00040703",
   341 => x"74200000",
   342 => x"787c5454",
   343 => x"7f7f0000",
   344 => x"387c4444",
   345 => x"7c380000",
   346 => x"00444444",
   347 => x"7c380000",
   348 => x"7f7f4444",
   349 => x"7c380000",
   350 => x"185c5454",
   351 => x"7e040000",
   352 => x"0005057f",
   353 => x"bc180000",
   354 => x"7cfca4a4",
   355 => x"7f7f0000",
   356 => x"787c0404",
   357 => x"00000000",
   358 => x"00407d3d",
   359 => x"80800000",
   360 => x"007dfd80",
   361 => x"7f7f0000",
   362 => x"446c3810",
   363 => x"00000000",
   364 => x"00407f3f",
   365 => x"0c7c7c00",
   366 => x"787c0c18",
   367 => x"7c7c0000",
   368 => x"787c0404",
   369 => x"7c380000",
   370 => x"387c4444",
   371 => x"fcfc0000",
   372 => x"183c2424",
   373 => x"3c180000",
   374 => x"fcfc2424",
   375 => x"7c7c0000",
   376 => x"080c0404",
   377 => x"5c480000",
   378 => x"20745454",
   379 => x"3f040000",
   380 => x"0044447f",
   381 => x"7c3c0000",
   382 => x"7c7c4040",
   383 => x"3c1c0000",
   384 => x"1c3c6060",
   385 => x"607c3c00",
   386 => x"3c7c6030",
   387 => x"386c4400",
   388 => x"446c3810",
   389 => x"bc1c0000",
   390 => x"1c3c60e0",
   391 => x"64440000",
   392 => x"444c5c74",
   393 => x"08080000",
   394 => x"4141773e",
   395 => x"00000000",
   396 => x"00007f7f",
   397 => x"41410000",
   398 => x"08083e77",
   399 => x"01010200",
   400 => x"01020203",
   401 => x"7f7f7f00",
   402 => x"7f7f7f7f",
   403 => x"1c080800",
   404 => x"7f3e3e1c",
   405 => x"3e7f7f7f",
   406 => x"081c1c3e",
   407 => x"18100008",
   408 => x"10187c7c",
   409 => x"30100000",
   410 => x"10307c7c",
   411 => x"60301000",
   412 => x"061e7860",
   413 => x"3c664200",
   414 => x"42663c18",
   415 => x"6a387800",
   416 => x"386cc6c2",
   417 => x"00006000",
   418 => x"60000060",
   419 => x"5b5e0e00",
   420 => x"1e0e5d5c",
   421 => x"c7c34c71",
   422 => x"c04dbfdf",
   423 => x"741ec04b",
   424 => x"87c702ab",
   425 => x"c048a6c4",
   426 => x"c487c578",
   427 => x"78c148a6",
   428 => x"731e66c4",
   429 => x"87dfee49",
   430 => x"e0c086c8",
   431 => x"87efef49",
   432 => x"6a4aa5c4",
   433 => x"87f0f049",
   434 => x"cb87c6f1",
   435 => x"c883c185",
   436 => x"ff04abb7",
   437 => x"262687c7",
   438 => x"264c264d",
   439 => x"1e4f264b",
   440 => x"c7c34a71",
   441 => x"c7c35ae3",
   442 => x"78c748e3",
   443 => x"87ddfe49",
   444 => x"731e4f26",
   445 => x"c04a711e",
   446 => x"d303aab7",
   447 => x"d1e9c287",
   448 => x"87c405bf",
   449 => x"87c24bc1",
   450 => x"e9c24bc0",
   451 => x"87c45bd5",
   452 => x"5ad5e9c2",
   453 => x"bfd1e9c2",
   454 => x"c19ac14a",
   455 => x"ec49a2c0",
   456 => x"48fc87e8",
   457 => x"bfd1e9c2",
   458 => x"87effe78",
   459 => x"c44a711e",
   460 => x"49721e66",
   461 => x"2687e2e6",
   462 => x"c21e4f26",
   463 => x"49bfd1e9",
   464 => x"87f2daff",
   465 => x"48d7c7c3",
   466 => x"c378bfe8",
   467 => x"ec48d3c7",
   468 => x"c7c378bf",
   469 => x"494abfd7",
   470 => x"c899ffc3",
   471 => x"48722ab7",
   472 => x"c7c3b071",
   473 => x"4f2658df",
   474 => x"5c5b5e0e",
   475 => x"4b710e5d",
   476 => x"c387c7ff",
   477 => x"c048d2c7",
   478 => x"ff497350",
   479 => x"7087d7da",
   480 => x"9cc24c49",
   481 => x"cb49eecb",
   482 => x"497087cf",
   483 => x"d2c7c34d",
   484 => x"c105bf97",
   485 => x"66d087e4",
   486 => x"dbc7c349",
   487 => x"d70599bf",
   488 => x"4966d487",
   489 => x"bfd3c7c3",
   490 => x"87cc0599",
   491 => x"d9ff4973",
   492 => x"987087e4",
   493 => x"87c2c102",
   494 => x"fdfd4cc1",
   495 => x"ca497587",
   496 => x"987087e3",
   497 => x"c387c602",
   498 => x"c148d2c7",
   499 => x"d2c7c350",
   500 => x"c005bf97",
   501 => x"c7c387e4",
   502 => x"d049bfdb",
   503 => x"ff059966",
   504 => x"c7c387d6",
   505 => x"d449bfd3",
   506 => x"ff059966",
   507 => x"497387ca",
   508 => x"87e2d8ff",
   509 => x"fe059870",
   510 => x"487487fe",
   511 => x"0e87d8fb",
   512 => x"5d5c5b5e",
   513 => x"c086f40e",
   514 => x"bfec4c4d",
   515 => x"48a6c47e",
   516 => x"bfdfc7c3",
   517 => x"c01ec178",
   518 => x"fd49c71e",
   519 => x"86c887ca",
   520 => x"ce029870",
   521 => x"fb49ff87",
   522 => x"dac187c8",
   523 => x"e5d7ff49",
   524 => x"c34dc187",
   525 => x"bf97d2c7",
   526 => x"d087c302",
   527 => x"c7c387c5",
   528 => x"c24bbfd7",
   529 => x"05bfd1e9",
   530 => x"c387ebc0",
   531 => x"d7ff49fd",
   532 => x"fac387c4",
   533 => x"fdd6ff49",
   534 => x"c3497387",
   535 => x"1e7199ff",
   536 => x"c7fb49c0",
   537 => x"c8497387",
   538 => x"1e7129b7",
   539 => x"fbfa49c1",
   540 => x"c686c887",
   541 => x"c7c387c1",
   542 => x"9b4bbfdb",
   543 => x"c287dd02",
   544 => x"49bfcde9",
   545 => x"7087dec7",
   546 => x"87c40598",
   547 => x"87d24bc0",
   548 => x"c749e0c2",
   549 => x"e9c287c3",
   550 => x"87c658d1",
   551 => x"48cde9c2",
   552 => x"497378c0",
   553 => x"ce0599c2",
   554 => x"49ebc387",
   555 => x"87e6d5ff",
   556 => x"99c24970",
   557 => x"fb87c202",
   558 => x"c149734c",
   559 => x"87ce0599",
   560 => x"ff49f4c3",
   561 => x"7087cfd5",
   562 => x"0299c249",
   563 => x"4cfa87c2",
   564 => x"99c84973",
   565 => x"c387ce05",
   566 => x"d4ff49f5",
   567 => x"497087f8",
   568 => x"d50299c2",
   569 => x"e3c7c387",
   570 => x"87ca02bf",
   571 => x"c388c148",
   572 => x"c058e7c7",
   573 => x"4cff87c2",
   574 => x"49734dc1",
   575 => x"ce0599c4",
   576 => x"49f2c387",
   577 => x"87ced4ff",
   578 => x"99c24970",
   579 => x"c387dc02",
   580 => x"7ebfe3c7",
   581 => x"a8b7c748",
   582 => x"87cbc003",
   583 => x"80c1486e",
   584 => x"58e7c7c3",
   585 => x"fe87c2c0",
   586 => x"c34dc14c",
   587 => x"d3ff49fd",
   588 => x"497087e4",
   589 => x"c00299c2",
   590 => x"c7c387d5",
   591 => x"c002bfe3",
   592 => x"c7c387c9",
   593 => x"78c048e3",
   594 => x"fd87c2c0",
   595 => x"c34dc14c",
   596 => x"d3ff49fa",
   597 => x"497087c0",
   598 => x"c00299c2",
   599 => x"c7c387d9",
   600 => x"c748bfe3",
   601 => x"c003a8b7",
   602 => x"c7c387c9",
   603 => x"78c748e3",
   604 => x"fc87c2c0",
   605 => x"c04dc14c",
   606 => x"c003acb7",
   607 => x"66c487d1",
   608 => x"82d8c14a",
   609 => x"c6c0026a",
   610 => x"744b6a87",
   611 => x"c00f7349",
   612 => x"1ef0c31e",
   613 => x"f749dac1",
   614 => x"86c887ce",
   615 => x"c0029870",
   616 => x"a6c887e2",
   617 => x"e3c7c348",
   618 => x"66c878bf",
   619 => x"c491cb49",
   620 => x"80714866",
   621 => x"bf6e7e70",
   622 => x"87c8c002",
   623 => x"c84bbf6e",
   624 => x"0f734966",
   625 => x"c0029d75",
   626 => x"c7c387c8",
   627 => x"f249bfe3",
   628 => x"e9c287fb",
   629 => x"c002bfd5",
   630 => x"c24987dd",
   631 => x"987087c7",
   632 => x"87d3c002",
   633 => x"bfe3c7c3",
   634 => x"87e1f249",
   635 => x"c1f449c0",
   636 => x"d5e9c287",
   637 => x"f478c048",
   638 => x"87dbf38e",
   639 => x"5c5b5e0e",
   640 => x"711e0e5d",
   641 => x"dfc7c34c",
   642 => x"cdc149bf",
   643 => x"d1c14da1",
   644 => x"747e6981",
   645 => x"87cf029c",
   646 => x"744ba5c4",
   647 => x"dfc7c37b",
   648 => x"faf249bf",
   649 => x"747b6e87",
   650 => x"87c4059c",
   651 => x"87c24bc0",
   652 => x"49734bc1",
   653 => x"d487fbf2",
   654 => x"87c70266",
   655 => x"7087da49",
   656 => x"c087c24a",
   657 => x"d9e9c24a",
   658 => x"caf2265a",
   659 => x"00000087",
   660 => x"00000000",
   661 => x"00000000",
   662 => x"4a711e00",
   663 => x"49bfc8ff",
   664 => x"2648a172",
   665 => x"c8ff1e4f",
   666 => x"c0fe89bf",
   667 => x"c0c0c0c0",
   668 => x"87c401a9",
   669 => x"87c24ac0",
   670 => x"48724ac1",
   671 => x"5e0e4f26",
   672 => x"0e5d5c5b",
   673 => x"d4ff4b71",
   674 => x"4866d04c",
   675 => x"49d678c0",
   676 => x"87cbd8ff",
   677 => x"6c7cffc3",
   678 => x"99ffc349",
   679 => x"c3494d71",
   680 => x"e0c199f0",
   681 => x"87cb05a9",
   682 => x"6c7cffc3",
   683 => x"d098c348",
   684 => x"c3780866",
   685 => x"4a6c7cff",
   686 => x"c331c849",
   687 => x"4a6c7cff",
   688 => x"4972b271",
   689 => x"ffc331c8",
   690 => x"714a6c7c",
   691 => x"c84972b2",
   692 => x"7cffc331",
   693 => x"b2714a6c",
   694 => x"c048d0ff",
   695 => x"9b7378e0",
   696 => x"7287c202",
   697 => x"2648757b",
   698 => x"264c264d",
   699 => x"1e4f264b",
   700 => x"5e0e4f26",
   701 => x"f80e5c5b",
   702 => x"c81e7686",
   703 => x"fdfd49a6",
   704 => x"7086c487",
   705 => x"c2486e4b",
   706 => x"f0c203a8",
   707 => x"c34a7387",
   708 => x"d0c19af0",
   709 => x"87c702aa",
   710 => x"05aae0c1",
   711 => x"7387dec2",
   712 => x"0299c849",
   713 => x"c6ff87c3",
   714 => x"c34c7387",
   715 => x"05acc29c",
   716 => x"c487c2c1",
   717 => x"31c94966",
   718 => x"66c41e71",
   719 => x"c392d44a",
   720 => x"7249e7c7",
   721 => x"d7fafd81",
   722 => x"ff49d887",
   723 => x"c887d0d5",
   724 => x"f5c21ec0",
   725 => x"d6fd49de",
   726 => x"d0ff87d2",
   727 => x"78e0c048",
   728 => x"1edef5c2",
   729 => x"d44a66cc",
   730 => x"e7c7c392",
   731 => x"fd817249",
   732 => x"cc87def8",
   733 => x"05acc186",
   734 => x"c487c2c1",
   735 => x"31c94966",
   736 => x"66c41e71",
   737 => x"c392d44a",
   738 => x"7249e7c7",
   739 => x"cff9fd81",
   740 => x"def5c287",
   741 => x"4a66c81e",
   742 => x"c7c392d4",
   743 => x"817249e7",
   744 => x"87def6fd",
   745 => x"d3ff49d7",
   746 => x"c0c887f5",
   747 => x"def5c21e",
   748 => x"d0d4fd49",
   749 => x"ff86cc87",
   750 => x"e0c048d0",
   751 => x"fc8ef878",
   752 => x"5e0e87e7",
   753 => x"0e5d5c5b",
   754 => x"ff4d711e",
   755 => x"66d44cd4",
   756 => x"b7c3487e",
   757 => x"87c506a8",
   758 => x"e2c148c0",
   759 => x"fe497587",
   760 => x"7587e3c7",
   761 => x"4b66c41e",
   762 => x"c7c393d4",
   763 => x"497383e7",
   764 => x"87f9f1fd",
   765 => x"4b6b83c8",
   766 => x"c848d0ff",
   767 => x"7cdd78e1",
   768 => x"ffc34973",
   769 => x"737c7199",
   770 => x"29b7c849",
   771 => x"7199ffc3",
   772 => x"d049737c",
   773 => x"ffc329b7",
   774 => x"737c7199",
   775 => x"29b7d849",
   776 => x"7cc07c71",
   777 => x"7c7c7c7c",
   778 => x"7c7c7c7c",
   779 => x"c07c7c7c",
   780 => x"66c478e0",
   781 => x"ff49dc1e",
   782 => x"c887c9d2",
   783 => x"26487386",
   784 => x"1e87e4fa",
   785 => x"bff4f4c2",
   786 => x"c2b9c149",
   787 => x"ff59f8f4",
   788 => x"ffc348d4",
   789 => x"48d0ff78",
   790 => x"ff78e1c8",
   791 => x"78c148d4",
   792 => x"787131c4",
   793 => x"c048d0ff",
   794 => x"4f2678e0",
   795 => x"c5f2c21e",
   796 => x"d4c2c31e",
   797 => x"f4effd49",
   798 => x"7086c487",
   799 => x"87c30298",
   800 => x"2687c0ff",
   801 => x"4b35314f",
   802 => x"20205a48",
   803 => x"47464320",
   804 => x"4a711e00",
   805 => x"c349a2c4",
   806 => x"6a48fac6",
   807 => x"c1496978",
   808 => x"f8f4c2b9",
   809 => x"87dbfe59",
   810 => x"87cad1ff",
   811 => x"4f2648c1",
   812 => x"c44a711e",
   813 => x"c6c349a2",
   814 => x"c27abffa",
   815 => x"79bff4f4",
   816 => x"711e4f26",
   817 => x"c0029a4a",
   818 => x"c31e87ec",
   819 => x"fd49d4c2",
   820 => x"c487daee",
   821 => x"02987086",
   822 => x"f5c287dc",
   823 => x"c2c31ede",
   824 => x"f1fd49d4",
   825 => x"86c487dc",
   826 => x"c9029870",
   827 => x"def5c287",
   828 => x"87ddfe49",
   829 => x"48c087c2",
   830 => x"711e4f26",
   831 => x"c0029a4a",
   832 => x"c31e87ee",
   833 => x"fd49d4c2",
   834 => x"c487e2ed",
   835 => x"02987086",
   836 => x"f5c287de",
   837 => x"d7fe49de",
   838 => x"def5c287",
   839 => x"d4c2c31e",
   840 => x"ecf1fd49",
   841 => x"7086c487",
   842 => x"87c40298",
   843 => x"87c248c1",
   844 => x"4f2648c0",
   845 => x"00000000",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
