library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.demistify_config_pkg.all;

-- -----------------------------------------------------------------------

entity de0nano_top is
	port
	(
		CLOCK_50		: IN STD_LOGIC;
		KEY			: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		SW				: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		LED			: OUT STD_LOGIC_VECTOR(7 DOWNTO 0) := (others=>'0');

		DRAM_CLK		: OUT STD_LOGIC;
		DRAM_CKE		: OUT STD_LOGIC;
		DRAM_ADDR	: OUT STD_LOGIC_VECTOR(12 DOWNTO 0);
		DRAM_BA		: OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		DRAM_DQ		: INOUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		DRAM_LDQM	: OUT STD_LOGIC;
		DRAM_UDQM	: OUT STD_LOGIC;
		DRAM_CS_N	: OUT STD_LOGIC;
		DRAM_WE_N	: OUT STD_LOGIC;
		DRAM_CAS_N	: OUT STD_LOGIC;
		DRAM_RAS_N	: OUT STD_LOGIC;
		
--		EPCS_DATA0	: INOUT std_logic_vector;
--		EPCS_DCLK	: INOUT std_logic_vector;
--		EPCS_NVCSO	: OUT std_logic_vector;
--		EPCS_ASDO	: OUT std_logic_vector;

		I2C_SCLK		: OUT STD_LOGIC;
		I2C_SDAT		: INOUT STD_LOGIC;

		G_SENSOR_INT: IN STD_LOGIC;
		G_SENSOR_CS_N: OUT STD_LOGIC;
		
		ADC_CS_N		: IN STD_LOGIC;
		ADC_SADDR	: OUT STD_LOGIC;
		ADC_SCLK		: OUT STD_LOGIC;
		ADC_SDAT		: IN STD_LOGIC;

		GPIO_0		: INOUT STD_LOGIC_VECTOR(33 DOWNTO 0) := (others => 'Z');
		GPIO_1		: INOUT STD_LOGIC_VECTOR(33 DOWNTO 0) := (others => 'Z');
		GPIO_2		: INOUT STD_LOGIC_VECTOR(12 DOWNTO 0) := (others => 'Z');
		GPIO_0_IN	: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		GPIO_1_IN	: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		GPIO_2_IN	: IN STD_LOGIC_VECTOR(2 DOWNTO 0)
	);
END entity;

architecture RTL of de0nano_top is
   constant reset_cycles : integer := 131071;
	
-- System clocks

	signal locked : std_logic;
	signal reset_n : std_logic;

--	signal slowclk : std_logic;
--	signal fastclk : std_logic;
--	signal pll_locked : std_logic;

-- SPI signals

	signal sd_clk : std_logic;
	signal sd_cs : std_logic;
	signal sd_mosi : std_logic;
	signal sd_miso : std_logic;
	
-- internal SPI signals
	
	signal spi_do : std_logic;
	signal spi_toguest : std_logic;
	signal spi_fromguest : std_logic;
	signal spi_ss2 : std_logic;
	signal spi_ss3 : std_logic;
	signal spi_ss4 : std_logic;
	signal conf_data0 : std_logic;
	signal spi_clk_int : std_logic;

-- PS/2 Keyboard socket - used for second mouse
	alias ps2_keyboard_clk : std_logic is GPIO_1(29); -- Dar
	alias ps2_keyboard_dat : std_logic is GPIO_1(27); -- Dar

	signal ps2_keyboard_clk_in : std_logic;
	signal ps2_keyboard_dat_in : std_logic;
	signal ps2_keyboard_clk_out : std_logic;
	signal ps2_keyboard_dat_out : std_logic;

-- PS/2 Mouse
	alias ps2_mouse_clk : std_logic is GPIO_1(33); -- Dar
	alias ps2_mouse_dat : std_logic is GPIO_1(31); -- Dar

	signal ps2_mouse_clk_in: std_logic;
	signal ps2_mouse_dat_in: std_logic;
	signal ps2_mouse_clk_out: std_logic;
	signal ps2_mouse_dat_out: std_logic;

	signal intercept : std_logic;
	
-- Video
	signal vga_red: std_logic_vector(7 downto 0);
	signal vga_green: std_logic_vector(7 downto 0);
	signal vga_blue: std_logic_vector(7 downto 0);
	signal vga_hsync : std_logic;
	signal vga_vsync : std_logic;

-- RS232 serial
	signal rs232_rxd : std_logic;
	signal rs232_txd : std_logic;

	signal sigma_l : std_logic;
	signal sigma_r : std_logic;
	
-- IO

	signal joya : std_logic_vector(7 downto 0);
	signal joyb : std_logic_vector(7 downto 0);
	signal joyc : std_logic_vector(7 downto 0);
	signal joyd : std_logic_vector(7 downto 0);

	signal uart_rxd : std_logic;
	signal uart_txd : std_logic;

	COMPONENT throbber
		PORT
		(
			clk		:	 IN STD_LOGIC;
			reset_n		:	 IN STD_LOGIC;
			q		:	 OUT STD_LOGIC
		);
	END COMPONENT;
	signal act_led : std_logic;

begin

--JOYSTICK
joya <= "111" & GPIO_1_IN(1) & GPIO_1_IN(0) & GPIO_1(6) & GPIO_1(8) & GPIO_1(10);     -- Dar
joyb <= "111" & GPIO_1(12) & GPIO_1(14) & GPIO_1(16) & GPIO_1(18) & GPIO_1(20); -- Dar

-- AUDIO
GPIO_1(2) <= sigma_l; -- Dar
GPIO_1(4) <= sigma_l; -- Dar

-- SPI
GPIO_1(28)<=sd_cs;   -- Dar
GPIO_1(26)<=sd_mosi; -- Dar
GPIO_1(24)<='Z';     -- Dar
sd_miso<=GPIO_1(24); -- Dar
GPIO_1(32)<=sd_clk;  -- Dar

-- PCXT serial
--GPIO_1(20) <= uart_txd;  -- Dar
--GPIO_1(21) <= 'Z';       -- Dar
--uart_rxd <= GPIO_1(21);  -- Dar

-- MCU serial
GPIO_0(2) <= rs232_txd;
GPIO_0(3) <= 'Z';
rs232_rxd <= GPIO_0(3);


--GPIO_1(22) <= uart_rts;  -- Dar
--GPIO_1(23) <= 'Z';       -- Dar
--uart_cts <= GPIO_1(23);  -- Dar

-- External devices tied to GPIOs

ps2_mouse_dat_in<=ps2_mouse_dat;
ps2_mouse_dat <= '0' when ps2_mouse_dat_out='0' else 'Z';
ps2_mouse_clk_in<=ps2_mouse_clk;
ps2_mouse_clk <= '0' when ps2_mouse_clk_out='0' else 'Z';

ps2_keyboard_dat_in<=ps2_keyboard_dat;
ps2_keyboard_dat <= '0' when ps2_keyboard_dat_out='0' else 'Z';
ps2_keyboard_clk_in<=ps2_keyboard_clk;
ps2_keyboard_clk <= '0' when ps2_keyboard_clk_out='0' else 'Z';

GPIO_1(25) <= vga_red(7); -- Dar
GPIO_1(23) <= vga_red(6); -- Dar
GPIO_1(21) <= vga_red(5); -- Dar
GPIO_1(19) <= vga_red(4); -- Dar
GPIO_1(17) <= vga_green(7); -- Dar
GPIO_1(15) <= vga_green(6); -- Dar
GPIO_1(13) <= vga_green(5); -- Dar
GPIO_1(11) <= vga_green(4); -- Dar
GPIO_1(9) <= vga_blue(7); -- Dar
GPIO_1(7) <= vga_blue(6); -- Dar
GPIO_1(5) <= vga_blue(5); -- Dar
GPIO_1(3) <= vga_blue(4); -- Dar
GPIO_1(1)<=vga_hsync;								-- Dar
GPIO_1(0)<=vga_vsync;								-- Dar


-- Generate clocks

guest: entity work.c64_mist
	PORT map
	(
--		CLOCK_27 => CLOCK_50&CLOCK_50, -- Comment out one of these lines to match the guest core.
		CLOCK_27 => CLOCK_50,
--		RESET_N => reset_n,
		LED => LED(0),
		-- clocks
		SDRAM_DQ => DRAM_DQ,
		SDRAM_A => DRAM_ADDR,
		SDRAM_DQML => DRAM_LDQM,
		SDRAM_DQMH => DRAM_UDQM,
		SDRAM_nWE => DRAM_WE_N,
		SDRAM_nCAS => DRAM_CAS_N,
		SDRAM_nRAS => DRAM_RAS_N,
		SDRAM_nCS => DRAM_CS_N,
		SDRAM_BA => DRAM_BA,
		SDRAM_CLK => DRAM_CLK,
		SDRAM_CKE => DRAM_CKE,
		
		SPI_DO => spi_do,
		SPI_DI => spi_toguest,
		SPI_SCK => spi_clk_int,
		SPI_SS2	=> spi_ss2,
		SPI_SS3 => spi_ss3,
		SPI_SS4 => spi_ss4,
		
		CONF_DATA0 => conf_data0,

		VGA_HS => vga_hsync,
		VGA_VS => vga_vsync,
		VGA_R => vga_red(7 downto 2),
		VGA_G => vga_green(7 downto 2),
		VGA_B => vga_blue(7 downto 2),
		AUDIO_L => sigma_l,
		AUDIO_R => sigma_r,
		
		UART_RX => '0',
		UART_TX => open
--		PS2K_CLK => ps2_keyboard_clk_in or intercept, -- Block keyboard when OSD is active
--		PS2K_DAT => ps2_keyboard_dat_in,
--		PS2M_CLK => ps2_mouse_clk_in,
--		PS2M_DAT => ps2_mouse_dat_in
);

-- Pass internal signals to external SPI interface
sd_clk <= spi_clk_int;
spi_do <= sd_miso when spi_ss4='0' else 'Z';
spi_fromguest <= spi_do;

controller : entity work.substitute_mcu
	generic map (
		sysclk_frequency => 500,
		--		SPI_FASTBIT=>3,
		--		SPI_INTERNALBIT=>2,		--keyb beeps if I discomment these two lines
		debug     => false,
		jtag_uart => false
	)
	port map (
		clk => CLOCK_50,
		reset_in => KEY(0),
		reset_out => reset_n,

		-- SPI signals
		spi_miso => sd_miso,
		spi_mosi	=> sd_mosi,
		spi_clk => spi_clk_int,
		spi_cs => sd_cs,
		spi_fromguest => spi_fromguest,
		spi_toguest => spi_toguest,
		spi_ss2 => spi_ss2,
		spi_ss3 => spi_ss3,
		spi_ss4 => spi_ss4,
		conf_data0 => conf_data0,
		
		-- PS/2 signals
		ps2k_clk_in => ps2_keyboard_clk_in,
		ps2k_dat_in => ps2_keyboard_dat_in,
		ps2k_clk_out => ps2_keyboard_clk_out,
		ps2k_dat_out => ps2_keyboard_dat_out,
		ps2m_clk_in => ps2_mouse_clk_in,
		ps2m_dat_in => ps2_mouse_dat_in,
		ps2m_clk_out => ps2_mouse_clk_out,
		ps2m_dat_out => ps2_mouse_dat_out,

		joy1 => joya,
		joy2 => joyb,
		buttons => (0=>KEY(1),others=>'1'),

		-- UART
		rxd => rs232_rxd,
		txd => rs232_txd,
		intercept => intercept
);

I2C_SCLK			<= '0';
I2C_SDAT			<= 'Z';
G_SENSOR_CS_N	<= '1';
ADC_SADDR		<= '0';
ADC_SCLK			<= '0';

end rtl;

