
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"71",x"78",x"c1",x"48"),
     1 => (x"c6",x"c0",x"02",x"99"),
     2 => (x"4c",x"f2",x"c0",x"87"),
     3 => (x"d7",x"87",x"c3",x"c0"),
     4 => (x"49",x"74",x"4c",x"dc"),
     5 => (x"87",x"c1",x"e9",x"c0"),
     6 => (x"c6",x"c3",x"49",x"70"),
     7 => (x"db",x"c1",x"59",x"fa"),
     8 => (x"e2",x"c6",x"c3",x"87"),
     9 => (x"87",x"de",x"ee",x"49"),
    10 => (x"02",x"9b",x"4b",x"70"),
    11 => (x"c2",x"87",x"ee",x"c0"),
    12 => (x"b7",x"bf",x"cb",x"c2"),
    13 => (x"e4",x"c0",x"03",x"ab"),
    14 => (x"f6",x"c6",x"c3",x"87"),
    15 => (x"e8",x"c0",x"49",x"bf"),
    16 => (x"98",x"70",x"87",x"e3"),
    17 => (x"87",x"f4",x"c0",x"02"),
    18 => (x"c2",x"c2",x"48",x"c7"),
    19 => (x"c2",x"88",x"bf",x"cb"),
    20 => (x"c3",x"58",x"cf",x"c2"),
    21 => (x"e9",x"49",x"e2",x"c6"),
    22 => (x"df",x"c0",x"87",x"df"),
    23 => (x"49",x"dc",x"d7",x"87"),
    24 => (x"87",x"f5",x"e7",x"c0"),
    25 => (x"c6",x"c3",x"49",x"70"),
    26 => (x"c2",x"c2",x"59",x"fa"),
    27 => (x"b7",x"4a",x"bf",x"cb"),
    28 => (x"c7",x"c0",x"04",x"ab"),
    29 => (x"d5",x"f8",x"49",x"87"),
    30 => (x"87",x"e5",x"fe",x"87"),
    31 => (x"00",x"87",x"dd",x"f9"),
    32 => (x"00",x"00",x"00",x"00"),
    33 => (x"00",x"00",x"00",x"00"),
    34 => (x"04",x"00",x"00",x"00"),
    35 => (x"01",x"00",x"00",x"00"),
    36 => (x"f3",x"08",x"82",x"ff"),
    37 => (x"f3",x"64",x"f3",x"c8"),
    38 => (x"81",x"01",x"f2",x"50"),
    39 => (x"1e",x"00",x"f4",x"01"),
    40 => (x"c8",x"48",x"d0",x"ff"),
    41 => (x"48",x"71",x"78",x"e1"),
    42 => (x"78",x"08",x"d4",x"ff"),
    43 => (x"ff",x"1e",x"4f",x"26"),
    44 => (x"e1",x"c8",x"48",x"d0"),
    45 => (x"ff",x"48",x"71",x"78"),
    46 => (x"c4",x"78",x"08",x"d4"),
    47 => (x"d4",x"ff",x"48",x"66"),
    48 => (x"4f",x"26",x"78",x"08"),
    49 => (x"c4",x"4a",x"71",x"1e"),
    50 => (x"72",x"1e",x"49",x"66"),
    51 => (x"87",x"de",x"ff",x"49"),
    52 => (x"c0",x"48",x"d0",x"ff"),
    53 => (x"26",x"26",x"78",x"e0"),
    54 => (x"1e",x"73",x"1e",x"4f"),
    55 => (x"66",x"c8",x"4b",x"71"),
    56 => (x"4a",x"73",x"1e",x"49"),
    57 => (x"49",x"a2",x"e0",x"c1"),
    58 => (x"26",x"87",x"d9",x"ff"),
    59 => (x"4d",x"26",x"87",x"c4"),
    60 => (x"4b",x"26",x"4c",x"26"),
    61 => (x"ff",x"1e",x"4f",x"26"),
    62 => (x"ff",x"c3",x"4a",x"d4"),
    63 => (x"48",x"d0",x"ff",x"7a"),
    64 => (x"de",x"78",x"e1",x"c8"),
    65 => (x"fa",x"c6",x"c3",x"7a"),
    66 => (x"48",x"49",x"7a",x"bf"),
    67 => (x"7a",x"70",x"28",x"c8"),
    68 => (x"28",x"d0",x"48",x"71"),
    69 => (x"48",x"71",x"7a",x"70"),
    70 => (x"7a",x"70",x"28",x"d8"),
    71 => (x"bf",x"fe",x"c6",x"c3"),
    72 => (x"c8",x"48",x"49",x"7a"),
    73 => (x"71",x"7a",x"70",x"28"),
    74 => (x"70",x"28",x"d0",x"48"),
    75 => (x"d8",x"48",x"71",x"7a"),
    76 => (x"ff",x"7a",x"70",x"28"),
    77 => (x"e0",x"c0",x"48",x"d0"),
    78 => (x"1e",x"4f",x"26",x"78"),
    79 => (x"4a",x"71",x"1e",x"73"),
    80 => (x"bf",x"fa",x"c6",x"c3"),
    81 => (x"c0",x"2b",x"72",x"4b"),
    82 => (x"ce",x"04",x"aa",x"e0"),
    83 => (x"c0",x"49",x"72",x"87"),
    84 => (x"c6",x"c3",x"89",x"e0"),
    85 => (x"71",x"4b",x"bf",x"fe"),
    86 => (x"c0",x"87",x"cf",x"2b"),
    87 => (x"89",x"72",x"49",x"e0"),
    88 => (x"bf",x"fe",x"c6",x"c3"),
    89 => (x"70",x"30",x"71",x"48"),
    90 => (x"66",x"c8",x"b3",x"49"),
    91 => (x"c4",x"48",x"73",x"9b"),
    92 => (x"26",x"4d",x"26",x"87"),
    93 => (x"26",x"4b",x"26",x"4c"),
    94 => (x"5b",x"5e",x"0e",x"4f"),
    95 => (x"ec",x"0e",x"5d",x"5c"),
    96 => (x"c3",x"4b",x"71",x"86"),
    97 => (x"7e",x"bf",x"fa",x"c6"),
    98 => (x"c0",x"2c",x"73",x"4c"),
    99 => (x"c0",x"04",x"ab",x"e0"),
   100 => (x"a6",x"c4",x"87",x"e0"),
   101 => (x"73",x"78",x"c0",x"48"),
   102 => (x"89",x"e0",x"c0",x"49"),
   103 => (x"e4",x"c0",x"4a",x"71"),
   104 => (x"30",x"72",x"48",x"66"),
   105 => (x"c3",x"58",x"a6",x"cc"),
   106 => (x"4d",x"bf",x"fe",x"c6"),
   107 => (x"c0",x"2c",x"71",x"4c"),
   108 => (x"49",x"73",x"87",x"e4"),
   109 => (x"48",x"66",x"e4",x"c0"),
   110 => (x"a6",x"c8",x"30",x"71"),
   111 => (x"49",x"e0",x"c0",x"58"),
   112 => (x"e4",x"c0",x"89",x"73"),
   113 => (x"28",x"71",x"48",x"66"),
   114 => (x"c3",x"58",x"a6",x"cc"),
   115 => (x"4d",x"bf",x"fe",x"c6"),
   116 => (x"70",x"30",x"71",x"48"),
   117 => (x"e4",x"c0",x"b4",x"49"),
   118 => (x"84",x"c1",x"9c",x"66"),
   119 => (x"ac",x"66",x"e8",x"c0"),
   120 => (x"c0",x"87",x"c2",x"04"),
   121 => (x"ab",x"e0",x"c0",x"4c"),
   122 => (x"cc",x"87",x"d3",x"04"),
   123 => (x"78",x"c0",x"48",x"a6"),
   124 => (x"e0",x"c0",x"49",x"73"),
   125 => (x"71",x"48",x"74",x"89"),
   126 => (x"58",x"a6",x"d4",x"30"),
   127 => (x"49",x"73",x"87",x"d5"),
   128 => (x"30",x"71",x"48",x"74"),
   129 => (x"c0",x"58",x"a6",x"d0"),
   130 => (x"89",x"73",x"49",x"e0"),
   131 => (x"28",x"71",x"48",x"74"),
   132 => (x"c4",x"58",x"a6",x"d4"),
   133 => (x"ba",x"ff",x"4a",x"66"),
   134 => (x"66",x"c8",x"9a",x"6e"),
   135 => (x"75",x"b9",x"ff",x"49"),
   136 => (x"cc",x"48",x"72",x"99"),
   137 => (x"c6",x"c3",x"b0",x"66"),
   138 => (x"48",x"71",x"58",x"fe"),
   139 => (x"c3",x"b0",x"66",x"d0"),
   140 => (x"fb",x"58",x"c2",x"c7"),
   141 => (x"8e",x"ec",x"87",x"c0"),
   142 => (x"1e",x"87",x"f6",x"fc"),
   143 => (x"c8",x"48",x"d0",x"ff"),
   144 => (x"48",x"71",x"78",x"c9"),
   145 => (x"78",x"08",x"d4",x"ff"),
   146 => (x"71",x"1e",x"4f",x"26"),
   147 => (x"87",x"eb",x"49",x"4a"),
   148 => (x"c8",x"48",x"d0",x"ff"),
   149 => (x"1e",x"4f",x"26",x"78"),
   150 => (x"4b",x"71",x"1e",x"73"),
   151 => (x"bf",x"ce",x"c7",x"c3"),
   152 => (x"c2",x"87",x"c3",x"02"),
   153 => (x"d0",x"ff",x"87",x"eb"),
   154 => (x"78",x"c9",x"c8",x"48"),
   155 => (x"e0",x"c0",x"49",x"73"),
   156 => (x"48",x"d4",x"ff",x"b1"),
   157 => (x"c7",x"c3",x"78",x"71"),
   158 => (x"78",x"c0",x"48",x"c2"),
   159 => (x"c5",x"02",x"66",x"c8"),
   160 => (x"49",x"ff",x"c3",x"87"),
   161 => (x"49",x"c0",x"87",x"c2"),
   162 => (x"59",x"ca",x"c7",x"c3"),
   163 => (x"c6",x"02",x"66",x"cc"),
   164 => (x"d5",x"d5",x"c5",x"87"),
   165 => (x"cf",x"87",x"c4",x"4a"),
   166 => (x"c3",x"4a",x"ff",x"ff"),
   167 => (x"c3",x"5a",x"ce",x"c7"),
   168 => (x"c1",x"48",x"ce",x"c7"),
   169 => (x"26",x"87",x"c4",x"78"),
   170 => (x"26",x"4c",x"26",x"4d"),
   171 => (x"0e",x"4f",x"26",x"4b"),
   172 => (x"5d",x"5c",x"5b",x"5e"),
   173 => (x"c3",x"4a",x"71",x"0e"),
   174 => (x"4c",x"bf",x"ca",x"c7"),
   175 => (x"cb",x"02",x"9a",x"72"),
   176 => (x"91",x"c8",x"49",x"87"),
   177 => (x"4b",x"cd",x"c9",x"c2"),
   178 => (x"87",x"c4",x"83",x"71"),
   179 => (x"4b",x"cd",x"cd",x"c2"),
   180 => (x"49",x"13",x"4d",x"c0"),
   181 => (x"c7",x"c3",x"99",x"74"),
   182 => (x"ff",x"b9",x"bf",x"c6"),
   183 => (x"78",x"71",x"48",x"d4"),
   184 => (x"85",x"2c",x"b7",x"c1"),
   185 => (x"04",x"ad",x"b7",x"c8"),
   186 => (x"c7",x"c3",x"87",x"e8"),
   187 => (x"c8",x"48",x"bf",x"c2"),
   188 => (x"c6",x"c7",x"c3",x"80"),
   189 => (x"87",x"ef",x"fe",x"58"),
   190 => (x"71",x"1e",x"73",x"1e"),
   191 => (x"9a",x"4a",x"13",x"4b"),
   192 => (x"72",x"87",x"cb",x"02"),
   193 => (x"87",x"e7",x"fe",x"49"),
   194 => (x"05",x"9a",x"4a",x"13"),
   195 => (x"da",x"fe",x"87",x"f5"),
   196 => (x"c7",x"c3",x"1e",x"87"),
   197 => (x"c3",x"49",x"bf",x"c2"),
   198 => (x"c1",x"48",x"c2",x"c7"),
   199 => (x"c0",x"c4",x"78",x"a1"),
   200 => (x"db",x"03",x"a9",x"b7"),
   201 => (x"48",x"d4",x"ff",x"87"),
   202 => (x"bf",x"c6",x"c7",x"c3"),
   203 => (x"c2",x"c7",x"c3",x"78"),
   204 => (x"c7",x"c3",x"49",x"bf"),
   205 => (x"a1",x"c1",x"48",x"c2"),
   206 => (x"b7",x"c0",x"c4",x"78"),
   207 => (x"87",x"e5",x"04",x"a9"),
   208 => (x"c8",x"48",x"d0",x"ff"),
   209 => (x"ce",x"c7",x"c3",x"78"),
   210 => (x"26",x"78",x"c0",x"48"),
   211 => (x"00",x"00",x"00",x"4f"),
   212 => (x"00",x"00",x"00",x"00"),
   213 => (x"00",x"00",x"00",x"00"),
   214 => (x"00",x"00",x"5f",x"5f"),
   215 => (x"03",x"03",x"00",x"00"),
   216 => (x"00",x"03",x"03",x"00"),
   217 => (x"7f",x"7f",x"14",x"00"),
   218 => (x"14",x"7f",x"7f",x"14"),
   219 => (x"2e",x"24",x"00",x"00"),
   220 => (x"12",x"3a",x"6b",x"6b"),
   221 => (x"36",x"6a",x"4c",x"00"),
   222 => (x"32",x"56",x"6c",x"18"),
   223 => (x"4f",x"7e",x"30",x"00"),
   224 => (x"68",x"3a",x"77",x"59"),
   225 => (x"04",x"00",x"00",x"40"),
   226 => (x"00",x"00",x"03",x"07"),
   227 => (x"1c",x"00",x"00",x"00"),
   228 => (x"00",x"41",x"63",x"3e"),
   229 => (x"41",x"00",x"00",x"00"),
   230 => (x"00",x"1c",x"3e",x"63"),
   231 => (x"3e",x"2a",x"08",x"00"),
   232 => (x"2a",x"3e",x"1c",x"1c"),
   233 => (x"08",x"08",x"00",x"08"),
   234 => (x"08",x"08",x"3e",x"3e"),
   235 => (x"80",x"00",x"00",x"00"),
   236 => (x"00",x"00",x"60",x"e0"),
   237 => (x"08",x"08",x"00",x"00"),
   238 => (x"08",x"08",x"08",x"08"),
   239 => (x"00",x"00",x"00",x"00"),
   240 => (x"00",x"00",x"60",x"60"),
   241 => (x"30",x"60",x"40",x"00"),
   242 => (x"03",x"06",x"0c",x"18"),
   243 => (x"7f",x"3e",x"00",x"01"),
   244 => (x"3e",x"7f",x"4d",x"59"),
   245 => (x"06",x"04",x"00",x"00"),
   246 => (x"00",x"00",x"7f",x"7f"),
   247 => (x"63",x"42",x"00",x"00"),
   248 => (x"46",x"4f",x"59",x"71"),
   249 => (x"63",x"22",x"00",x"00"),
   250 => (x"36",x"7f",x"49",x"49"),
   251 => (x"16",x"1c",x"18",x"00"),
   252 => (x"10",x"7f",x"7f",x"13"),
   253 => (x"67",x"27",x"00",x"00"),
   254 => (x"39",x"7d",x"45",x"45"),
   255 => (x"7e",x"3c",x"00",x"00"),
   256 => (x"30",x"79",x"49",x"4b"),
   257 => (x"01",x"01",x"00",x"00"),
   258 => (x"07",x"0f",x"79",x"71"),
   259 => (x"7f",x"36",x"00",x"00"),
   260 => (x"36",x"7f",x"49",x"49"),
   261 => (x"4f",x"06",x"00",x"00"),
   262 => (x"1e",x"3f",x"69",x"49"),
   263 => (x"00",x"00",x"00",x"00"),
   264 => (x"00",x"00",x"66",x"66"),
   265 => (x"80",x"00",x"00",x"00"),
   266 => (x"00",x"00",x"66",x"e6"),
   267 => (x"08",x"08",x"00",x"00"),
   268 => (x"22",x"22",x"14",x"14"),
   269 => (x"14",x"14",x"00",x"00"),
   270 => (x"14",x"14",x"14",x"14"),
   271 => (x"22",x"22",x"00",x"00"),
   272 => (x"08",x"08",x"14",x"14"),
   273 => (x"03",x"02",x"00",x"00"),
   274 => (x"06",x"0f",x"59",x"51"),
   275 => (x"41",x"7f",x"3e",x"00"),
   276 => (x"1e",x"1f",x"55",x"5d"),
   277 => (x"7f",x"7e",x"00",x"00"),
   278 => (x"7e",x"7f",x"09",x"09"),
   279 => (x"7f",x"7f",x"00",x"00"),
   280 => (x"36",x"7f",x"49",x"49"),
   281 => (x"3e",x"1c",x"00",x"00"),
   282 => (x"41",x"41",x"41",x"63"),
   283 => (x"7f",x"7f",x"00",x"00"),
   284 => (x"1c",x"3e",x"63",x"41"),
   285 => (x"7f",x"7f",x"00",x"00"),
   286 => (x"41",x"41",x"49",x"49"),
   287 => (x"7f",x"7f",x"00",x"00"),
   288 => (x"01",x"01",x"09",x"09"),
   289 => (x"7f",x"3e",x"00",x"00"),
   290 => (x"7a",x"7b",x"49",x"41"),
   291 => (x"7f",x"7f",x"00",x"00"),
   292 => (x"7f",x"7f",x"08",x"08"),
   293 => (x"41",x"00",x"00",x"00"),
   294 => (x"00",x"41",x"7f",x"7f"),
   295 => (x"60",x"20",x"00",x"00"),
   296 => (x"3f",x"7f",x"40",x"40"),
   297 => (x"08",x"7f",x"7f",x"00"),
   298 => (x"41",x"63",x"36",x"1c"),
   299 => (x"7f",x"7f",x"00",x"00"),
   300 => (x"40",x"40",x"40",x"40"),
   301 => (x"06",x"7f",x"7f",x"00"),
   302 => (x"7f",x"7f",x"06",x"0c"),
   303 => (x"06",x"7f",x"7f",x"00"),
   304 => (x"7f",x"7f",x"18",x"0c"),
   305 => (x"7f",x"3e",x"00",x"00"),
   306 => (x"3e",x"7f",x"41",x"41"),
   307 => (x"7f",x"7f",x"00",x"00"),
   308 => (x"06",x"0f",x"09",x"09"),
   309 => (x"41",x"7f",x"3e",x"00"),
   310 => (x"40",x"7e",x"7f",x"61"),
   311 => (x"7f",x"7f",x"00",x"00"),
   312 => (x"66",x"7f",x"19",x"09"),
   313 => (x"6f",x"26",x"00",x"00"),
   314 => (x"32",x"7b",x"59",x"4d"),
   315 => (x"01",x"01",x"00",x"00"),
   316 => (x"01",x"01",x"7f",x"7f"),
   317 => (x"7f",x"3f",x"00",x"00"),
   318 => (x"3f",x"7f",x"40",x"40"),
   319 => (x"3f",x"0f",x"00",x"00"),
   320 => (x"0f",x"3f",x"70",x"70"),
   321 => (x"30",x"7f",x"7f",x"00"),
   322 => (x"7f",x"7f",x"30",x"18"),
   323 => (x"36",x"63",x"41",x"00"),
   324 => (x"63",x"36",x"1c",x"1c"),
   325 => (x"06",x"03",x"01",x"41"),
   326 => (x"03",x"06",x"7c",x"7c"),
   327 => (x"59",x"71",x"61",x"01"),
   328 => (x"41",x"43",x"47",x"4d"),
   329 => (x"7f",x"00",x"00",x"00"),
   330 => (x"00",x"41",x"41",x"7f"),
   331 => (x"06",x"03",x"01",x"00"),
   332 => (x"60",x"30",x"18",x"0c"),
   333 => (x"41",x"00",x"00",x"40"),
   334 => (x"00",x"7f",x"7f",x"41"),
   335 => (x"06",x"0c",x"08",x"00"),
   336 => (x"08",x"0c",x"06",x"03"),
   337 => (x"80",x"80",x"80",x"00"),
   338 => (x"80",x"80",x"80",x"80"),
   339 => (x"00",x"00",x"00",x"00"),
   340 => (x"00",x"04",x"07",x"03"),
   341 => (x"74",x"20",x"00",x"00"),
   342 => (x"78",x"7c",x"54",x"54"),
   343 => (x"7f",x"7f",x"00",x"00"),
   344 => (x"38",x"7c",x"44",x"44"),
   345 => (x"7c",x"38",x"00",x"00"),
   346 => (x"00",x"44",x"44",x"44"),
   347 => (x"7c",x"38",x"00",x"00"),
   348 => (x"7f",x"7f",x"44",x"44"),
   349 => (x"7c",x"38",x"00",x"00"),
   350 => (x"18",x"5c",x"54",x"54"),
   351 => (x"7e",x"04",x"00",x"00"),
   352 => (x"00",x"05",x"05",x"7f"),
   353 => (x"bc",x"18",x"00",x"00"),
   354 => (x"7c",x"fc",x"a4",x"a4"),
   355 => (x"7f",x"7f",x"00",x"00"),
   356 => (x"78",x"7c",x"04",x"04"),
   357 => (x"00",x"00",x"00",x"00"),
   358 => (x"00",x"40",x"7d",x"3d"),
   359 => (x"80",x"80",x"00",x"00"),
   360 => (x"00",x"7d",x"fd",x"80"),
   361 => (x"7f",x"7f",x"00",x"00"),
   362 => (x"44",x"6c",x"38",x"10"),
   363 => (x"00",x"00",x"00",x"00"),
   364 => (x"00",x"40",x"7f",x"3f"),
   365 => (x"0c",x"7c",x"7c",x"00"),
   366 => (x"78",x"7c",x"0c",x"18"),
   367 => (x"7c",x"7c",x"00",x"00"),
   368 => (x"78",x"7c",x"04",x"04"),
   369 => (x"7c",x"38",x"00",x"00"),
   370 => (x"38",x"7c",x"44",x"44"),
   371 => (x"fc",x"fc",x"00",x"00"),
   372 => (x"18",x"3c",x"24",x"24"),
   373 => (x"3c",x"18",x"00",x"00"),
   374 => (x"fc",x"fc",x"24",x"24"),
   375 => (x"7c",x"7c",x"00",x"00"),
   376 => (x"08",x"0c",x"04",x"04"),
   377 => (x"5c",x"48",x"00",x"00"),
   378 => (x"20",x"74",x"54",x"54"),
   379 => (x"3f",x"04",x"00",x"00"),
   380 => (x"00",x"44",x"44",x"7f"),
   381 => (x"7c",x"3c",x"00",x"00"),
   382 => (x"7c",x"7c",x"40",x"40"),
   383 => (x"3c",x"1c",x"00",x"00"),
   384 => (x"1c",x"3c",x"60",x"60"),
   385 => (x"60",x"7c",x"3c",x"00"),
   386 => (x"3c",x"7c",x"60",x"30"),
   387 => (x"38",x"6c",x"44",x"00"),
   388 => (x"44",x"6c",x"38",x"10"),
   389 => (x"bc",x"1c",x"00",x"00"),
   390 => (x"1c",x"3c",x"60",x"e0"),
   391 => (x"64",x"44",x"00",x"00"),
   392 => (x"44",x"4c",x"5c",x"74"),
   393 => (x"08",x"08",x"00",x"00"),
   394 => (x"41",x"41",x"77",x"3e"),
   395 => (x"00",x"00",x"00",x"00"),
   396 => (x"00",x"00",x"7f",x"7f"),
   397 => (x"41",x"41",x"00",x"00"),
   398 => (x"08",x"08",x"3e",x"77"),
   399 => (x"01",x"01",x"02",x"00"),
   400 => (x"01",x"02",x"02",x"03"),
   401 => (x"7f",x"7f",x"7f",x"00"),
   402 => (x"7f",x"7f",x"7f",x"7f"),
   403 => (x"1c",x"08",x"08",x"00"),
   404 => (x"7f",x"3e",x"3e",x"1c"),
   405 => (x"3e",x"7f",x"7f",x"7f"),
   406 => (x"08",x"1c",x"1c",x"3e"),
   407 => (x"18",x"10",x"00",x"08"),
   408 => (x"10",x"18",x"7c",x"7c"),
   409 => (x"30",x"10",x"00",x"00"),
   410 => (x"10",x"30",x"7c",x"7c"),
   411 => (x"60",x"30",x"10",x"00"),
   412 => (x"06",x"1e",x"78",x"60"),
   413 => (x"3c",x"66",x"42",x"00"),
   414 => (x"42",x"66",x"3c",x"18"),
   415 => (x"6a",x"38",x"78",x"00"),
   416 => (x"38",x"6c",x"c6",x"c2"),
   417 => (x"00",x"00",x"60",x"00"),
   418 => (x"60",x"00",x"00",x"60"),
   419 => (x"5b",x"5e",x"0e",x"00"),
   420 => (x"1e",x"0e",x"5d",x"5c"),
   421 => (x"c7",x"c3",x"4c",x"71"),
   422 => (x"c0",x"4d",x"bf",x"df"),
   423 => (x"74",x"1e",x"c0",x"4b"),
   424 => (x"87",x"c7",x"02",x"ab"),
   425 => (x"c0",x"48",x"a6",x"c4"),
   426 => (x"c4",x"87",x"c5",x"78"),
   427 => (x"78",x"c1",x"48",x"a6"),
   428 => (x"73",x"1e",x"66",x"c4"),
   429 => (x"87",x"df",x"ee",x"49"),
   430 => (x"e0",x"c0",x"86",x"c8"),
   431 => (x"87",x"ef",x"ef",x"49"),
   432 => (x"6a",x"4a",x"a5",x"c4"),
   433 => (x"87",x"f0",x"f0",x"49"),
   434 => (x"cb",x"87",x"c6",x"f1"),
   435 => (x"c8",x"83",x"c1",x"85"),
   436 => (x"ff",x"04",x"ab",x"b7"),
   437 => (x"26",x"26",x"87",x"c7"),
   438 => (x"26",x"4c",x"26",x"4d"),
   439 => (x"1e",x"4f",x"26",x"4b"),
   440 => (x"c7",x"c3",x"4a",x"71"),
   441 => (x"c7",x"c3",x"5a",x"e3"),
   442 => (x"78",x"c7",x"48",x"e3"),
   443 => (x"87",x"dd",x"fe",x"49"),
   444 => (x"73",x"1e",x"4f",x"26"),
   445 => (x"c0",x"4a",x"71",x"1e"),
   446 => (x"d3",x"03",x"aa",x"b7"),
   447 => (x"d1",x"e9",x"c2",x"87"),
   448 => (x"87",x"c4",x"05",x"bf"),
   449 => (x"87",x"c2",x"4b",x"c1"),
   450 => (x"e9",x"c2",x"4b",x"c0"),
   451 => (x"87",x"c4",x"5b",x"d5"),
   452 => (x"5a",x"d5",x"e9",x"c2"),
   453 => (x"bf",x"d1",x"e9",x"c2"),
   454 => (x"c1",x"9a",x"c1",x"4a"),
   455 => (x"ec",x"49",x"a2",x"c0"),
   456 => (x"48",x"fc",x"87",x"e8"),
   457 => (x"bf",x"d1",x"e9",x"c2"),
   458 => (x"87",x"ef",x"fe",x"78"),
   459 => (x"c4",x"4a",x"71",x"1e"),
   460 => (x"49",x"72",x"1e",x"66"),
   461 => (x"26",x"87",x"e2",x"e6"),
   462 => (x"c2",x"1e",x"4f",x"26"),
   463 => (x"49",x"bf",x"d1",x"e9"),
   464 => (x"87",x"f2",x"da",x"ff"),
   465 => (x"48",x"d7",x"c7",x"c3"),
   466 => (x"c3",x"78",x"bf",x"e8"),
   467 => (x"ec",x"48",x"d3",x"c7"),
   468 => (x"c7",x"c3",x"78",x"bf"),
   469 => (x"49",x"4a",x"bf",x"d7"),
   470 => (x"c8",x"99",x"ff",x"c3"),
   471 => (x"48",x"72",x"2a",x"b7"),
   472 => (x"c7",x"c3",x"b0",x"71"),
   473 => (x"4f",x"26",x"58",x"df"),
   474 => (x"5c",x"5b",x"5e",x"0e"),
   475 => (x"4b",x"71",x"0e",x"5d"),
   476 => (x"c3",x"87",x"c7",x"ff"),
   477 => (x"c0",x"48",x"d2",x"c7"),
   478 => (x"ff",x"49",x"73",x"50"),
   479 => (x"70",x"87",x"d7",x"da"),
   480 => (x"9c",x"c2",x"4c",x"49"),
   481 => (x"cb",x"49",x"ee",x"cb"),
   482 => (x"49",x"70",x"87",x"cf"),
   483 => (x"d2",x"c7",x"c3",x"4d"),
   484 => (x"c1",x"05",x"bf",x"97"),
   485 => (x"66",x"d0",x"87",x"e4"),
   486 => (x"db",x"c7",x"c3",x"49"),
   487 => (x"d7",x"05",x"99",x"bf"),
   488 => (x"49",x"66",x"d4",x"87"),
   489 => (x"bf",x"d3",x"c7",x"c3"),
   490 => (x"87",x"cc",x"05",x"99"),
   491 => (x"d9",x"ff",x"49",x"73"),
   492 => (x"98",x"70",x"87",x"e4"),
   493 => (x"87",x"c2",x"c1",x"02"),
   494 => (x"fd",x"fd",x"4c",x"c1"),
   495 => (x"ca",x"49",x"75",x"87"),
   496 => (x"98",x"70",x"87",x"e3"),
   497 => (x"c3",x"87",x"c6",x"02"),
   498 => (x"c1",x"48",x"d2",x"c7"),
   499 => (x"d2",x"c7",x"c3",x"50"),
   500 => (x"c0",x"05",x"bf",x"97"),
   501 => (x"c7",x"c3",x"87",x"e4"),
   502 => (x"d0",x"49",x"bf",x"db"),
   503 => (x"ff",x"05",x"99",x"66"),
   504 => (x"c7",x"c3",x"87",x"d6"),
   505 => (x"d4",x"49",x"bf",x"d3"),
   506 => (x"ff",x"05",x"99",x"66"),
   507 => (x"49",x"73",x"87",x"ca"),
   508 => (x"87",x"e2",x"d8",x"ff"),
   509 => (x"fe",x"05",x"98",x"70"),
   510 => (x"48",x"74",x"87",x"fe"),
   511 => (x"0e",x"87",x"d8",x"fb"),
   512 => (x"5d",x"5c",x"5b",x"5e"),
   513 => (x"c0",x"86",x"f4",x"0e"),
   514 => (x"bf",x"ec",x"4c",x"4d"),
   515 => (x"48",x"a6",x"c4",x"7e"),
   516 => (x"bf",x"df",x"c7",x"c3"),
   517 => (x"c0",x"1e",x"c1",x"78"),
   518 => (x"fd",x"49",x"c7",x"1e"),
   519 => (x"86",x"c8",x"87",x"ca"),
   520 => (x"ce",x"02",x"98",x"70"),
   521 => (x"fb",x"49",x"ff",x"87"),
   522 => (x"da",x"c1",x"87",x"c8"),
   523 => (x"e5",x"d7",x"ff",x"49"),
   524 => (x"c3",x"4d",x"c1",x"87"),
   525 => (x"bf",x"97",x"d2",x"c7"),
   526 => (x"d0",x"87",x"c3",x"02"),
   527 => (x"c7",x"c3",x"87",x"c5"),
   528 => (x"c2",x"4b",x"bf",x"d7"),
   529 => (x"05",x"bf",x"d1",x"e9"),
   530 => (x"c3",x"87",x"eb",x"c0"),
   531 => (x"d7",x"ff",x"49",x"fd"),
   532 => (x"fa",x"c3",x"87",x"c4"),
   533 => (x"fd",x"d6",x"ff",x"49"),
   534 => (x"c3",x"49",x"73",x"87"),
   535 => (x"1e",x"71",x"99",x"ff"),
   536 => (x"c7",x"fb",x"49",x"c0"),
   537 => (x"c8",x"49",x"73",x"87"),
   538 => (x"1e",x"71",x"29",x"b7"),
   539 => (x"fb",x"fa",x"49",x"c1"),
   540 => (x"c6",x"86",x"c8",x"87"),
   541 => (x"c7",x"c3",x"87",x"c1"),
   542 => (x"9b",x"4b",x"bf",x"db"),
   543 => (x"c2",x"87",x"dd",x"02"),
   544 => (x"49",x"bf",x"cd",x"e9"),
   545 => (x"70",x"87",x"de",x"c7"),
   546 => (x"87",x"c4",x"05",x"98"),
   547 => (x"87",x"d2",x"4b",x"c0"),
   548 => (x"c7",x"49",x"e0",x"c2"),
   549 => (x"e9",x"c2",x"87",x"c3"),
   550 => (x"87",x"c6",x"58",x"d1"),
   551 => (x"48",x"cd",x"e9",x"c2"),
   552 => (x"49",x"73",x"78",x"c0"),
   553 => (x"ce",x"05",x"99",x"c2"),
   554 => (x"49",x"eb",x"c3",x"87"),
   555 => (x"87",x"e6",x"d5",x"ff"),
   556 => (x"99",x"c2",x"49",x"70"),
   557 => (x"fb",x"87",x"c2",x"02"),
   558 => (x"c1",x"49",x"73",x"4c"),
   559 => (x"87",x"ce",x"05",x"99"),
   560 => (x"ff",x"49",x"f4",x"c3"),
   561 => (x"70",x"87",x"cf",x"d5"),
   562 => (x"02",x"99",x"c2",x"49"),
   563 => (x"4c",x"fa",x"87",x"c2"),
   564 => (x"99",x"c8",x"49",x"73"),
   565 => (x"c3",x"87",x"ce",x"05"),
   566 => (x"d4",x"ff",x"49",x"f5"),
   567 => (x"49",x"70",x"87",x"f8"),
   568 => (x"d5",x"02",x"99",x"c2"),
   569 => (x"e3",x"c7",x"c3",x"87"),
   570 => (x"87",x"ca",x"02",x"bf"),
   571 => (x"c3",x"88",x"c1",x"48"),
   572 => (x"c0",x"58",x"e7",x"c7"),
   573 => (x"4c",x"ff",x"87",x"c2"),
   574 => (x"49",x"73",x"4d",x"c1"),
   575 => (x"ce",x"05",x"99",x"c4"),
   576 => (x"49",x"f2",x"c3",x"87"),
   577 => (x"87",x"ce",x"d4",x"ff"),
   578 => (x"99",x"c2",x"49",x"70"),
   579 => (x"c3",x"87",x"dc",x"02"),
   580 => (x"7e",x"bf",x"e3",x"c7"),
   581 => (x"a8",x"b7",x"c7",x"48"),
   582 => (x"87",x"cb",x"c0",x"03"),
   583 => (x"80",x"c1",x"48",x"6e"),
   584 => (x"58",x"e7",x"c7",x"c3"),
   585 => (x"fe",x"87",x"c2",x"c0"),
   586 => (x"c3",x"4d",x"c1",x"4c"),
   587 => (x"d3",x"ff",x"49",x"fd"),
   588 => (x"49",x"70",x"87",x"e4"),
   589 => (x"c0",x"02",x"99",x"c2"),
   590 => (x"c7",x"c3",x"87",x"d5"),
   591 => (x"c0",x"02",x"bf",x"e3"),
   592 => (x"c7",x"c3",x"87",x"c9"),
   593 => (x"78",x"c0",x"48",x"e3"),
   594 => (x"fd",x"87",x"c2",x"c0"),
   595 => (x"c3",x"4d",x"c1",x"4c"),
   596 => (x"d3",x"ff",x"49",x"fa"),
   597 => (x"49",x"70",x"87",x"c0"),
   598 => (x"c0",x"02",x"99",x"c2"),
   599 => (x"c7",x"c3",x"87",x"d9"),
   600 => (x"c7",x"48",x"bf",x"e3"),
   601 => (x"c0",x"03",x"a8",x"b7"),
   602 => (x"c7",x"c3",x"87",x"c9"),
   603 => (x"78",x"c7",x"48",x"e3"),
   604 => (x"fc",x"87",x"c2",x"c0"),
   605 => (x"c0",x"4d",x"c1",x"4c"),
   606 => (x"c0",x"03",x"ac",x"b7"),
   607 => (x"66",x"c4",x"87",x"d1"),
   608 => (x"82",x"d8",x"c1",x"4a"),
   609 => (x"c6",x"c0",x"02",x"6a"),
   610 => (x"74",x"4b",x"6a",x"87"),
   611 => (x"c0",x"0f",x"73",x"49"),
   612 => (x"1e",x"f0",x"c3",x"1e"),
   613 => (x"f7",x"49",x"da",x"c1"),
   614 => (x"86",x"c8",x"87",x"ce"),
   615 => (x"c0",x"02",x"98",x"70"),
   616 => (x"a6",x"c8",x"87",x"e2"),
   617 => (x"e3",x"c7",x"c3",x"48"),
   618 => (x"66",x"c8",x"78",x"bf"),
   619 => (x"c4",x"91",x"cb",x"49"),
   620 => (x"80",x"71",x"48",x"66"),
   621 => (x"bf",x"6e",x"7e",x"70"),
   622 => (x"87",x"c8",x"c0",x"02"),
   623 => (x"c8",x"4b",x"bf",x"6e"),
   624 => (x"0f",x"73",x"49",x"66"),
   625 => (x"c0",x"02",x"9d",x"75"),
   626 => (x"c7",x"c3",x"87",x"c8"),
   627 => (x"f2",x"49",x"bf",x"e3"),
   628 => (x"e9",x"c2",x"87",x"fb"),
   629 => (x"c0",x"02",x"bf",x"d5"),
   630 => (x"c2",x"49",x"87",x"dd"),
   631 => (x"98",x"70",x"87",x"c7"),
   632 => (x"87",x"d3",x"c0",x"02"),
   633 => (x"bf",x"e3",x"c7",x"c3"),
   634 => (x"87",x"e1",x"f2",x"49"),
   635 => (x"c1",x"f4",x"49",x"c0"),
   636 => (x"d5",x"e9",x"c2",x"87"),
   637 => (x"f4",x"78",x"c0",x"48"),
   638 => (x"87",x"db",x"f3",x"8e"),
   639 => (x"5c",x"5b",x"5e",x"0e"),
   640 => (x"71",x"1e",x"0e",x"5d"),
   641 => (x"df",x"c7",x"c3",x"4c"),
   642 => (x"cd",x"c1",x"49",x"bf"),
   643 => (x"d1",x"c1",x"4d",x"a1"),
   644 => (x"74",x"7e",x"69",x"81"),
   645 => (x"87",x"cf",x"02",x"9c"),
   646 => (x"74",x"4b",x"a5",x"c4"),
   647 => (x"df",x"c7",x"c3",x"7b"),
   648 => (x"fa",x"f2",x"49",x"bf"),
   649 => (x"74",x"7b",x"6e",x"87"),
   650 => (x"87",x"c4",x"05",x"9c"),
   651 => (x"87",x"c2",x"4b",x"c0"),
   652 => (x"49",x"73",x"4b",x"c1"),
   653 => (x"d4",x"87",x"fb",x"f2"),
   654 => (x"87",x"c7",x"02",x"66"),
   655 => (x"70",x"87",x"da",x"49"),
   656 => (x"c0",x"87",x"c2",x"4a"),
   657 => (x"d9",x"e9",x"c2",x"4a"),
   658 => (x"ca",x"f2",x"26",x"5a"),
   659 => (x"00",x"00",x"00",x"87"),
   660 => (x"00",x"00",x"00",x"00"),
   661 => (x"00",x"00",x"00",x"00"),
   662 => (x"4a",x"71",x"1e",x"00"),
   663 => (x"49",x"bf",x"c8",x"ff"),
   664 => (x"26",x"48",x"a1",x"72"),
   665 => (x"c8",x"ff",x"1e",x"4f"),
   666 => (x"c0",x"fe",x"89",x"bf"),
   667 => (x"c0",x"c0",x"c0",x"c0"),
   668 => (x"87",x"c4",x"01",x"a9"),
   669 => (x"87",x"c2",x"4a",x"c0"),
   670 => (x"48",x"72",x"4a",x"c1"),
   671 => (x"5e",x"0e",x"4f",x"26"),
   672 => (x"0e",x"5d",x"5c",x"5b"),
   673 => (x"d4",x"ff",x"4b",x"71"),
   674 => (x"48",x"66",x"d0",x"4c"),
   675 => (x"49",x"d6",x"78",x"c0"),
   676 => (x"87",x"cb",x"d8",x"ff"),
   677 => (x"6c",x"7c",x"ff",x"c3"),
   678 => (x"99",x"ff",x"c3",x"49"),
   679 => (x"c3",x"49",x"4d",x"71"),
   680 => (x"e0",x"c1",x"99",x"f0"),
   681 => (x"87",x"cb",x"05",x"a9"),
   682 => (x"6c",x"7c",x"ff",x"c3"),
   683 => (x"d0",x"98",x"c3",x"48"),
   684 => (x"c3",x"78",x"08",x"66"),
   685 => (x"4a",x"6c",x"7c",x"ff"),
   686 => (x"c3",x"31",x"c8",x"49"),
   687 => (x"4a",x"6c",x"7c",x"ff"),
   688 => (x"49",x"72",x"b2",x"71"),
   689 => (x"ff",x"c3",x"31",x"c8"),
   690 => (x"71",x"4a",x"6c",x"7c"),
   691 => (x"c8",x"49",x"72",x"b2"),
   692 => (x"7c",x"ff",x"c3",x"31"),
   693 => (x"b2",x"71",x"4a",x"6c"),
   694 => (x"c0",x"48",x"d0",x"ff"),
   695 => (x"9b",x"73",x"78",x"e0"),
   696 => (x"72",x"87",x"c2",x"02"),
   697 => (x"26",x"48",x"75",x"7b"),
   698 => (x"26",x"4c",x"26",x"4d"),
   699 => (x"1e",x"4f",x"26",x"4b"),
   700 => (x"5e",x"0e",x"4f",x"26"),
   701 => (x"f8",x"0e",x"5c",x"5b"),
   702 => (x"c8",x"1e",x"76",x"86"),
   703 => (x"fd",x"fd",x"49",x"a6"),
   704 => (x"70",x"86",x"c4",x"87"),
   705 => (x"c2",x"48",x"6e",x"4b"),
   706 => (x"f0",x"c2",x"03",x"a8"),
   707 => (x"c3",x"4a",x"73",x"87"),
   708 => (x"d0",x"c1",x"9a",x"f0"),
   709 => (x"87",x"c7",x"02",x"aa"),
   710 => (x"05",x"aa",x"e0",x"c1"),
   711 => (x"73",x"87",x"de",x"c2"),
   712 => (x"02",x"99",x"c8",x"49"),
   713 => (x"c6",x"ff",x"87",x"c3"),
   714 => (x"c3",x"4c",x"73",x"87"),
   715 => (x"05",x"ac",x"c2",x"9c"),
   716 => (x"c4",x"87",x"c2",x"c1"),
   717 => (x"31",x"c9",x"49",x"66"),
   718 => (x"66",x"c4",x"1e",x"71"),
   719 => (x"c3",x"92",x"d4",x"4a"),
   720 => (x"72",x"49",x"e7",x"c7"),
   721 => (x"d7",x"fa",x"fd",x"81"),
   722 => (x"ff",x"49",x"d8",x"87"),
   723 => (x"c8",x"87",x"d0",x"d5"),
   724 => (x"f5",x"c2",x"1e",x"c0"),
   725 => (x"d6",x"fd",x"49",x"de"),
   726 => (x"d0",x"ff",x"87",x"d2"),
   727 => (x"78",x"e0",x"c0",x"48"),
   728 => (x"1e",x"de",x"f5",x"c2"),
   729 => (x"d4",x"4a",x"66",x"cc"),
   730 => (x"e7",x"c7",x"c3",x"92"),
   731 => (x"fd",x"81",x"72",x"49"),
   732 => (x"cc",x"87",x"de",x"f8"),
   733 => (x"05",x"ac",x"c1",x"86"),
   734 => (x"c4",x"87",x"c2",x"c1"),
   735 => (x"31",x"c9",x"49",x"66"),
   736 => (x"66",x"c4",x"1e",x"71"),
   737 => (x"c3",x"92",x"d4",x"4a"),
   738 => (x"72",x"49",x"e7",x"c7"),
   739 => (x"cf",x"f9",x"fd",x"81"),
   740 => (x"de",x"f5",x"c2",x"87"),
   741 => (x"4a",x"66",x"c8",x"1e"),
   742 => (x"c7",x"c3",x"92",x"d4"),
   743 => (x"81",x"72",x"49",x"e7"),
   744 => (x"87",x"de",x"f6",x"fd"),
   745 => (x"d3",x"ff",x"49",x"d7"),
   746 => (x"c0",x"c8",x"87",x"f5"),
   747 => (x"de",x"f5",x"c2",x"1e"),
   748 => (x"d0",x"d4",x"fd",x"49"),
   749 => (x"ff",x"86",x"cc",x"87"),
   750 => (x"e0",x"c0",x"48",x"d0"),
   751 => (x"fc",x"8e",x"f8",x"78"),
   752 => (x"5e",x"0e",x"87",x"e7"),
   753 => (x"0e",x"5d",x"5c",x"5b"),
   754 => (x"ff",x"4d",x"71",x"1e"),
   755 => (x"66",x"d4",x"4c",x"d4"),
   756 => (x"b7",x"c3",x"48",x"7e"),
   757 => (x"87",x"c5",x"06",x"a8"),
   758 => (x"e2",x"c1",x"48",x"c0"),
   759 => (x"fe",x"49",x"75",x"87"),
   760 => (x"75",x"87",x"e3",x"c7"),
   761 => (x"4b",x"66",x"c4",x"1e"),
   762 => (x"c7",x"c3",x"93",x"d4"),
   763 => (x"49",x"73",x"83",x"e7"),
   764 => (x"87",x"f9",x"f1",x"fd"),
   765 => (x"4b",x"6b",x"83",x"c8"),
   766 => (x"c8",x"48",x"d0",x"ff"),
   767 => (x"7c",x"dd",x"78",x"e1"),
   768 => (x"ff",x"c3",x"49",x"73"),
   769 => (x"73",x"7c",x"71",x"99"),
   770 => (x"29",x"b7",x"c8",x"49"),
   771 => (x"71",x"99",x"ff",x"c3"),
   772 => (x"d0",x"49",x"73",x"7c"),
   773 => (x"ff",x"c3",x"29",x"b7"),
   774 => (x"73",x"7c",x"71",x"99"),
   775 => (x"29",x"b7",x"d8",x"49"),
   776 => (x"7c",x"c0",x"7c",x"71"),
   777 => (x"7c",x"7c",x"7c",x"7c"),
   778 => (x"7c",x"7c",x"7c",x"7c"),
   779 => (x"c0",x"7c",x"7c",x"7c"),
   780 => (x"66",x"c4",x"78",x"e0"),
   781 => (x"ff",x"49",x"dc",x"1e"),
   782 => (x"c8",x"87",x"c9",x"d2"),
   783 => (x"26",x"48",x"73",x"86"),
   784 => (x"1e",x"87",x"e4",x"fa"),
   785 => (x"bf",x"f4",x"f4",x"c2"),
   786 => (x"c2",x"b9",x"c1",x"49"),
   787 => (x"ff",x"59",x"f8",x"f4"),
   788 => (x"ff",x"c3",x"48",x"d4"),
   789 => (x"48",x"d0",x"ff",x"78"),
   790 => (x"ff",x"78",x"e1",x"c8"),
   791 => (x"78",x"c1",x"48",x"d4"),
   792 => (x"78",x"71",x"31",x"c4"),
   793 => (x"c0",x"48",x"d0",x"ff"),
   794 => (x"4f",x"26",x"78",x"e0"),
   795 => (x"c5",x"f2",x"c2",x"1e"),
   796 => (x"d4",x"c2",x"c3",x"1e"),
   797 => (x"f4",x"ef",x"fd",x"49"),
   798 => (x"70",x"86",x"c4",x"87"),
   799 => (x"87",x"c3",x"02",x"98"),
   800 => (x"26",x"87",x"c0",x"ff"),
   801 => (x"4b",x"35",x"31",x"4f"),
   802 => (x"20",x"20",x"5a",x"48"),
   803 => (x"47",x"46",x"43",x"20"),
   804 => (x"4a",x"71",x"1e",x"00"),
   805 => (x"c3",x"49",x"a2",x"c4"),
   806 => (x"6a",x"48",x"fa",x"c6"),
   807 => (x"c1",x"49",x"69",x"78"),
   808 => (x"f8",x"f4",x"c2",x"b9"),
   809 => (x"87",x"db",x"fe",x"59"),
   810 => (x"87",x"ca",x"d1",x"ff"),
   811 => (x"4f",x"26",x"48",x"c1"),
   812 => (x"c4",x"4a",x"71",x"1e"),
   813 => (x"c6",x"c3",x"49",x"a2"),
   814 => (x"c2",x"7a",x"bf",x"fa"),
   815 => (x"79",x"bf",x"f4",x"f4"),
   816 => (x"71",x"1e",x"4f",x"26"),
   817 => (x"c0",x"02",x"9a",x"4a"),
   818 => (x"c3",x"1e",x"87",x"ec"),
   819 => (x"fd",x"49",x"d4",x"c2"),
   820 => (x"c4",x"87",x"da",x"ee"),
   821 => (x"02",x"98",x"70",x"86"),
   822 => (x"f5",x"c2",x"87",x"dc"),
   823 => (x"c2",x"c3",x"1e",x"de"),
   824 => (x"f1",x"fd",x"49",x"d4"),
   825 => (x"86",x"c4",x"87",x"dc"),
   826 => (x"c9",x"02",x"98",x"70"),
   827 => (x"de",x"f5",x"c2",x"87"),
   828 => (x"87",x"dd",x"fe",x"49"),
   829 => (x"48",x"c0",x"87",x"c2"),
   830 => (x"71",x"1e",x"4f",x"26"),
   831 => (x"c0",x"02",x"9a",x"4a"),
   832 => (x"c3",x"1e",x"87",x"ee"),
   833 => (x"fd",x"49",x"d4",x"c2"),
   834 => (x"c4",x"87",x"e2",x"ed"),
   835 => (x"02",x"98",x"70",x"86"),
   836 => (x"f5",x"c2",x"87",x"de"),
   837 => (x"d7",x"fe",x"49",x"de"),
   838 => (x"de",x"f5",x"c2",x"87"),
   839 => (x"d4",x"c2",x"c3",x"1e"),
   840 => (x"ec",x"f1",x"fd",x"49"),
   841 => (x"70",x"86",x"c4",x"87"),
   842 => (x"87",x"c4",x"02",x"98"),
   843 => (x"87",x"c2",x"48",x"c1"),
   844 => (x"4f",x"26",x"48",x"c0"),
   845 => (x"00",x"00",x"00",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

